`ifndef config_vh_
`define config_vh_

`define VERSION_MAJOR 8'd0
`define VERSION_MINOR 8'd8

`define REV_3_BOARD 1

`define VARIANT_SUFFIX_1 8'd0;
`define VARIANT_SUFFIX_2 8'd0;
`define VARIANT_SUFFIX_3 8'd0;
`define VARIANT_SUFFIX_4 8'd0;

`define WITH_EXTENSIONS 1
`define WITH_RAM 1
`define WITH_64K 1
`define WITH_DVI 1
`define GEN_LUMA_CHROMA 1
`define CONFIGURABLE_LUMAS 1
`define CONFIGURABLE_RGB 1
`define HAVE_EEPROM 1
`define HAVE_FLASH 1
`define NEED_RGB 1
`define GEN_RGB 1
`define HIRES_MODES
`define HIRES_RESET
`define WITH_MATH

`endif // config_vh_
