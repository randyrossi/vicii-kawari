`ifndef config_vh_
`define config_vh_

`define VERSION_MAJOR 8'd0
`define VERSION_MINOR 8'd8

`define REV_4S_BOARD 1
`define NO_CLOCK_MUX 1
`define GEN_LUMA_CHROMA 1

`endif // config_vh_
