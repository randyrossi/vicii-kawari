// This file is part of the vicii-kawari distribution
// (https://github.com/randyrossi/vicii-kawari)
// Copyright (c) 2022 Randy Rossi.
// 
// This program is free software: you can redistribute it and/or modify  
// it under the terms of the GNU General Public License as published by  
// the Free Software Foundation, version 3.
//
// This program is distributed in the hope that it will be useful, but 
// WITHOUT ANY WARRANTY; without even the implied warranty of 
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the GNU 
// General Public License for more details.
//
// You should have received a copy of the GNU General Public License 
// along with this program. If not, see <http://www.gnu.org/licenses/>.

`include "common.vh"

// NOTE: We reproduce the offscreen white pixel at hvisible_start
// that the real VICII's produces.  You can't see it on CRTs but it
// will show up on upscalers. It can be removed by getting rid of
// the three raster_x == hvisible_start conditions below for luma,
// phase and amplitude.

// Rev 4+ boards have luma sink capabilities to properly
// sink most current during h/v sync periods. Rev 3 board
// couldn't do this and the sync period was too 'hot' but
// still worked on most monitors.
`ifndef REV_3_BOARD
`define HAVE_LUMA_SINK 1
`endif

// A module that produces a luma/chroma signals.
module comp_sync(
           input clk_dot4x,
           input clk_col16x,
           input [9:0] raster_x,
           input [8:0] raster_y,
`ifdef GEN_LUMA_CHROMA
           input white_line,
           input ntsc_50,
           //input pal_60,
`ifdef HAVE_LUMA_SINK
           output reg luma_sink,
`endif
           output [5:0] luma_out,
           output reg [5:0] chroma_out,
           input [5:0] lumareg_o, // from registers base on pixel_color3
           input [7:0] phasereg_o, // from registers base on pixel_color3
           input [3:0] amplitudereg_o, // from registers base on pixel_color3
`ifdef CONFIGURABLE_LUMAS
           input [5:0] blanking_level,
           input [3:0] burst_amplitude,
`endif
`endif
           input [1:0] chip
       );

reg [5:0] luma;
reg [9:0] hvisible_end;
//reg [9:0] hsync_start; // now always 10'd10
reg [9:0] hsync_end;
reg [9:0] hvisible_start;
reg [8:0] vvisible_end;
reg [8:0] vblank_start;
//reg [8:0] vblank_end;
reg [8:0] vvisible_start;
reg hSync;
reg vSync;
reg native_active;

`ifdef GEN_LUMA_CHROMA
`ifdef HAVE_LUMA_SINK
assign luma_out = ~luma;
`else
assign luma_out = luma;
`endif
`endif

always @(posedge clk_dot4x)
begin
    // NOTE hsync_start is hard coded to 10'd10 to save a register. If this ever
    // changes, serration.v and equalization.v must also change.
    hSync <= raster_x >= 10'd10 /* hsync_start */ && raster_x < hsync_end;
    vSync <= (raster_y >= vvisible_end && raster_y <= vvisible_start);
    native_active <= ~(
                      (raster_x >= hvisible_end | raster_x < hvisible_start) |
                      (
                          ((raster_y == vvisible_end & raster_x < hvisible_end) | raster_y > vvisible_end) &
                          ((raster_y == vvisible_start & raster_x <= hvisible_start) | raster_y < vvisible_start)
                      )
                  );
end

// NTSC: Each x is ~122.2 ns (.1222 us)
// PAL : Each x is ~126.8 ns (.1268 us)
`ifdef SIMULATOR_BOARD
always @(posedge clk_dot4x)
`else
always @(chip)
`endif
case(chip)
    `CHIP6567R8:
    begin
        // 520x263
        hvisible_end = 10'd510;
        //hsync_start = 10'd10;
        hsync_end = 10'd49;      // .0075H
        hvisible_start = 10'd90;
        vvisible_end = 9'd13;
        vblank_start = 9'd14; // visible_end +9'd1
        //vblank_end = 9'd22; // vblank_start + 9'd8;
        vvisible_start = 9'd23; // vblank_end + 9'd1;
    end
    `CHIP6567R56A:
    begin
        // 512x262
        hvisible_end = 10'd502;
        //hsync_start = 10'd10;
        hsync_end = 10'd48;       // .0075H
        hvisible_start = 10'd90;
        vvisible_end = 9'd13;
        vblank_start = 9'd14; // visible_end +9'd1
        //vblank_end = 9'd22; // vblank_start + 9'd8;
        vvisible_start = 9'd23; // vblank_end + 9'd1;
    end
    `CHIP6569R1, `CHIP6569R3:
    begin
        // 504x312
        hvisible_end = 10'd494;
        //hsync_start = 10'd10;
        hsync_end = 10'd48;       // .0075H
        hvisible_start =  10'd90;
        vvisible_end = 9'd300;
        vblank_start = 9'd301; // visible_end +9'd1
        //vblank_end = 9'd309; // vblank_start + 9'd8;
        vvisible_start = 9'd310; // vblank_end + 9'd1;
    end
endcase

// NTSC
// 2.69us = 2690 ns
// 3.579545 Mhz = 279.3 ns period
// 2690 / 279.3 = 9.6 (need only 9 cycles of color clock)
//
// PAL
// 2.97us = 2970 ns
// 4.43361875 Mhz = 225.5 ns period
// 2970 / 225.5 = 13.1 (need only 9 cycles of color clock)

// Compute Equalization pulses
wire EQ, SE;
EqualizationPulse ueqp1
                  (
                      .clk_dot4x(clk_dot4x),
                      .raster_x(raster_x),
                      .chip(chip),
                      .EQ(EQ)
                  );

// Compute Serration pulses
SerrationPulse usep1
               (
                   .clk_dot4x(clk_dot4x),
                   .raster_x(raster_x),
                   .chip(chip),
                   .SE(SE)
               );

`ifdef GEN_LUMA_CHROMA

// Luma level of white burst on first visible pixel
`define WHITE_BURST 6'h3b

// If configurable, use register value.
// Otherwise, hard coded values.
`ifdef CONFIGURABLE_LUMAS
`define BLANKING_LEVEL blanking_level
`else
`ifdef REV_3_BOARD
`define BLANKING_LEVEL 6'd12
`else
`define BLANKING_LEVEL (chip[0] ? 6'h08 : 6'h18)
`endif
`endif

always @(posedge clk_dot4x)
begin
    begin
        case(raster_y)
            vblank_start: begin
               luma <= ~EQ ? `BLANKING_LEVEL : 6'd0;
`ifdef HAVE_LUMA_SINK
               luma_sink <= EQ;
`endif
            end
            vblank_start+1: begin
               luma <= ~EQ ? `BLANKING_LEVEL : 6'd0;
`ifdef HAVE_LUMA_SINK
               luma_sink <= EQ;
`endif
            end
            vblank_start+2: begin
               luma <= ~EQ ? `BLANKING_LEVEL : 6'd0;
`ifdef HAVE_LUMA_SINK
               luma_sink <= EQ;
`endif
            end
            vblank_start+3: begin
               luma <= ~SE ? `BLANKING_LEVEL : 6'd0;
`ifdef HAVE_LUMA_SINK
               luma_sink <= SE;
`endif
            end
            vblank_start+4: begin
               luma <= ~SE ? `BLANKING_LEVEL : 6'd0;
`ifdef HAVE_LUMA_SINK
               luma_sink <= SE;
`endif
            end
            vblank_start+5: begin
               luma <= ~SE ? `BLANKING_LEVEL : 6'd0;
`ifdef HAVE_LUMA_SINK
               luma_sink <= SE;
`endif
            end
            vblank_start+6: begin
               luma <= ~EQ ? `BLANKING_LEVEL : 6'd0;
`ifdef HAVE_LUMA_SINK
               luma_sink <= EQ;
`endif
            end
            vblank_start+7: begin
               luma <= ~EQ ? `BLANKING_LEVEL : 6'd0;
`ifdef HAVE_LUMA_SINK
               luma_sink <= EQ;
`endif
            end
            vblank_start+8: begin
               luma <= ~EQ ? `BLANKING_LEVEL : 6'd0;
`ifdef HAVE_LUMA_SINK
               luma_sink <= EQ;
`endif
            end
            // This is visible start but it should be a blank line
            vblank_start+9: begin
               luma <= ~hSync ? `BLANKING_LEVEL : 6'd0;
`ifdef HAVE_LUMA_SINK
               luma_sink <= hSync;
`endif
            end
            default: begin
                luma <= ~hSync ? (~native_active ? `BLANKING_LEVEL : ((raster_x == hvisible_start && white_line) ? `WHITE_BURST : lumareg_o)) : 6'd0;
`ifdef HAVE_LUMA_SINK
                luma_sink <= hSync;
`endif
            end
        endcase
    end
end

// Phase counter forms the first 4 bits of the index into our
// sine table of 256 entries.  Hence, it takes 16 samples from
// the sine table for every period of our 16x color clock and
// produces a 1x color clock wave.  The wave phase can be shifted
// by applying a phase offset of 8 bits.  The amplitude is selected
// out of the sine wave table rom by prefixing the 8 bits with
// an additional 4 bits of amplitude.
reg [3:0] phaseCounter;
reg [8:0] prev_raster_y;
reg [3:0] amplitude2;
reg [3:0] amplitude3;
reg [3:0] amplitude4;

always @(posedge clk_col16x)
begin
    phaseCounter <= phaseCounter + 4'd1;
end

`define NO_MODULATION 4'b0000

`ifdef CONFIGURABLE_LUMAS
`define BURST_AMPLITUDE burst_amplitude_16
`else
`define BURST_AMPLITUDE 4'd12
`endif

// Make this hsync_end + 4 ticks
// !!! Keep this valid for hsync_end set below:
// 6567R8 = 49 + 4 = 53
// 6567R56A = 48 + 4 = 52
// 6569R* = 48 + 4 = 52
`define BURST_START (chip_1_16x == `CHIP6567R8 ? 10'd53 : 10'd52)

(* async_reg = "true" *) reg [8:0] raster_y_16_1;
(* async_reg = "true" *) reg [8:0] raster_y_16;
(* async_reg = "true" *) reg [9:0] raster_x_16_1;
(* async_reg = "true" *) reg [9:0] raster_x_16;
(* async_reg = "true" *) reg native_active_16_1;
(* async_reg = "true" *) reg native_active_16;
(* async_reg = "true" *) reg vSync_16_1;
(* async_reg = "true" *) reg vSync_16;

// Handle domain crossing for registers we need from dot4x in a co16x block.
always @(posedge clk_col16x) raster_y_16_1 <= raster_y;
always @(posedge clk_col16x) raster_y_16 <= raster_y_16_1;
always @(posedge clk_col16x) raster_x_16_1 <= raster_x;
always @(posedge clk_col16x) raster_x_16 <= raster_x_16_1;
always @(posedge clk_col16x) native_active_16_1 <= native_active;
always @(posedge clk_col16x) native_active_16 <= native_active_16_1;
always @(posedge clk_col16x) vSync_16_1 <= vSync;
always @(posedge clk_col16x) vSync_16 <= vSync_16_1;

reg [7:0] burstCount;
reg [7:0] sineWaveAddr;
reg [11:0] sineROMAddr;
reg in_burst;
reg need_burst;
wire oddline;
assign oddline = raster_y_16[0];

(* async_reg = "true" *) reg [9:0] hvisible_start_16_1;
(* async_reg = "true" *) reg [9:0] hvisible_start_16;
always @(posedge clk_col16x) hvisible_start_16_1 <= hvisible_start;
always @(posedge clk_col16x) hvisible_start_16 <= hvisible_start_16_1;

// Handle domain crossing from dot4x to col16x
(* async_reg = "true" *) reg [7:0] phasereg_o2;
(* async_reg = "true" *) reg [7:0] phasereg_16;
always @(posedge clk_col16x) phasereg_o2 <= phasereg_o;
always @(posedge clk_col16x) phasereg_16 <= (raster_x_16 == hvisible_start_16 && white_line_16) ? 8'h0 : phasereg_o2;

(* async_reg = "true" *) reg [3:0] amplitudereg_o2;
(* async_reg = "true" *) reg [3:0] amplitudereg_16;
always @(posedge clk_col16x) amplitudereg_o2 <=  amplitudereg_o;
always @(posedge clk_col16x) amplitudereg_16 <= (raster_x_16 == hvisible_start_16 && white_line_16) ? 4'h0 : amplitudereg_o2;

`ifdef CONFIGURABLE_LUMAS
(* async_reg = "true" *) reg [3:0] burst_amplitude_ms;
(* async_reg = "true" *) reg [3:0] burst_amplitude_16;
always @(posedge clk_col16x) burst_amplitude_ms <=  burst_amplitude;
always @(posedge clk_col16x) burst_amplitude_16 <= burst_amplitude_ms;
`endif

(* async_reg = "true" *) reg colsel_0;
(* async_reg = "true" *) reg colsel_1;
always @(posedge clk_col16x) colsel_0 <= chip[0] ? (~ntsc_50) : 1'b0; // was (pal_60);
always @(posedge clk_col16x) colsel_1 <= colsel_0;

(* async_reg = "true" *) reg[1:0] chip_0_16x;
(* async_reg = "true" *) reg[1:0] chip_1_16x;
always @(posedge clk_col16x) chip_0_16x <= chip;
always @(posedge clk_col16x) chip_1_16x <= chip_0_16x;

(* async_reg = "true" *) reg white_line_ms;
(* async_reg = "true" *) reg white_line_16;
always @(posedge clk_col16x) white_line_ms <= white_line;
always @(posedge clk_col16x) white_line_16 <= white_line_ms;

reg [8:0] chroma9;

always @(posedge clk_col16x)
begin
    if (raster_y_16 != prev_raster_y) begin
        need_burst <= 1;
    end
    prev_raster_y <= raster_y_16;

    if (raster_x_16 >= `BURST_START && need_burst)
        in_burst <= 1;

    if (in_burst)
    begin
        // This is supposed to be 9 periods according to video specs but the
        // original chip does more like 20. I noticed that if we only do 9 and
        // use the PAL clock from the motherboard, we produce a B/W image.
        // Increased to 15 periods for PAL
        // One less for NTSC
        if ((chip_1_16x[0] && burstCount == 240) || (~chip_1_16x[0] && burstCount == 224))
        begin
            in_burst <= 0;
            need_burst <= 0;
            burstCount <= 0;
        end else begin
            burstCount <= burstCount + 1'b1;
        end
    end

    // Use amplitude from table lookup inside active region.  For burst, use
    // 4'b0100. Otherwise, amplitude should be 4'b0000 representing no
    // modulation.
    amplitude2 = vSync_16 ?
               `NO_MODULATION :
               (native_active_16 ?
                amplitudereg_16 :
                (in_burst ? `BURST_AMPLITUDE : `NO_MODULATION));

    amplitude3 <= amplitude2;
    amplitude4 <= amplitude3;
    // Figure out the entry within one of the sine wave tables.
    // For NTSC: Burst phase is always 180 degrees (128 offset)
    // For PAL: Burst phase alternates between 135 and -135 (96 & 160 offsets).
    /* verilator lint_off WIDTH */
    sineWaveAddr = {phaseCounter, 4'b0} +
                 (
                     native_active_16 ?
                     (colsel_1 ?
                      (oddline ? 8'd255 - phasereg_16 :  phasereg_16) : /* pal */
                      phasereg_16) :                                    /* ntsc */
                     (colsel_1 ?
                      (oddline ? 8'd160 : 8'd96) :                      /* pal */
                      8'd128                                            /* ntsc */
                     )
                 );

    /* verilator lint_on WIDTH */
    // Prefix with amplitude selector. This is our ROM address.
    sineROMAddr <= {amplitude2, sineWaveAddr };

    // Chroma is centered at 32 for no amplitude. (top 6 bits of 256 offset)
    // Make the decision to output chroma or zero level baseed on the amplitude that
    // was used to determine the chroma9 lookup (which was two ticks ago, one tick to set
    // the address and another to get the data)
    chroma_out <= (amplitude4 == `NO_MODULATION) ? 6'd32 : chroma9[8:3];
end

// Retrieve wave value from addr calculated from amplitude, phaseCounter and
// phaseOffset.
always @(sineROMAddr)
begin
    case (sineROMAddr)
        12'd0: chroma9 = 9'b000000000;
        12'd1: chroma9 = 9'b000000000;
        12'd2: chroma9 = 9'b000000000;
        12'd3: chroma9 = 9'b000000000;
        12'd4: chroma9 = 9'b000000000;
        12'd5: chroma9 = 9'b000000000;
        12'd6: chroma9 = 9'b000000000;
        12'd7: chroma9 = 9'b000000000;
        12'd8: chroma9 = 9'b000000000;
        12'd9: chroma9 = 9'b000000000;
        12'd10: chroma9 = 9'b000000000;
        12'd11: chroma9 = 9'b000000000;
        12'd12: chroma9 = 9'b000000000;
        12'd13: chroma9 = 9'b000000000;
        12'd14: chroma9 = 9'b000000000;
        12'd15: chroma9 = 9'b000000000;
        12'd16: chroma9 = 9'b000000000;
        12'd17: chroma9 = 9'b000000000;
        12'd18: chroma9 = 9'b000000000;
        12'd19: chroma9 = 9'b000000000;
        12'd20: chroma9 = 9'b000000000;
        12'd21: chroma9 = 9'b000000000;
        12'd22: chroma9 = 9'b000000000;
        12'd23: chroma9 = 9'b000000000;
        12'd24: chroma9 = 9'b000000000;
        12'd25: chroma9 = 9'b000000000;
        12'd26: chroma9 = 9'b000000000;
        12'd27: chroma9 = 9'b000000000;
        12'd28: chroma9 = 9'b000000000;
        12'd29: chroma9 = 9'b000000000;
        12'd30: chroma9 = 9'b000000000;
        12'd31: chroma9 = 9'b000000000;
        12'd32: chroma9 = 9'b000000000;
        12'd33: chroma9 = 9'b000000000;
        12'd34: chroma9 = 9'b000000000;
        12'd35: chroma9 = 9'b000000000;
        12'd36: chroma9 = 9'b000000000;
        12'd37: chroma9 = 9'b000000000;
        12'd38: chroma9 = 9'b000000000;
        12'd39: chroma9 = 9'b000000000;
        12'd40: chroma9 = 9'b000000000;
        12'd41: chroma9 = 9'b000000000;
        12'd42: chroma9 = 9'b000000000;
        12'd43: chroma9 = 9'b000000000;
        12'd44: chroma9 = 9'b000000000;
        12'd45: chroma9 = 9'b000000000;
        12'd46: chroma9 = 9'b000000000;
        12'd47: chroma9 = 9'b000000000;
        12'd48: chroma9 = 9'b000000000;
        12'd49: chroma9 = 9'b000000000;
        12'd50: chroma9 = 9'b000000000;
        12'd51: chroma9 = 9'b000000000;
        12'd52: chroma9 = 9'b000000000;
        12'd53: chroma9 = 9'b000000000;
        12'd54: chroma9 = 9'b000000000;
        12'd55: chroma9 = 9'b000000000;
        12'd56: chroma9 = 9'b000000000;
        12'd57: chroma9 = 9'b000000000;
        12'd58: chroma9 = 9'b000000000;
        12'd59: chroma9 = 9'b000000000;
        12'd60: chroma9 = 9'b000000000;
        12'd61: chroma9 = 9'b000000000;
        12'd62: chroma9 = 9'b000000000;
        12'd63: chroma9 = 9'b000000000;
        12'd64: chroma9 = 9'b000000000;
        12'd65: chroma9 = 9'b000000000;
        12'd66: chroma9 = 9'b000000000;
        12'd67: chroma9 = 9'b000000000;
        12'd68: chroma9 = 9'b000000000;
        12'd69: chroma9 = 9'b000000000;
        12'd70: chroma9 = 9'b000000000;
        12'd71: chroma9 = 9'b000000000;
        12'd72: chroma9 = 9'b000000000;
        12'd73: chroma9 = 9'b000000000;
        12'd74: chroma9 = 9'b000000000;
        12'd75: chroma9 = 9'b000000000;
        12'd76: chroma9 = 9'b000000000;
        12'd77: chroma9 = 9'b000000000;
        12'd78: chroma9 = 9'b000000000;
        12'd79: chroma9 = 9'b000000000;
        12'd80: chroma9 = 9'b000000000;
        12'd81: chroma9 = 9'b000000000;
        12'd82: chroma9 = 9'b000000000;
        12'd83: chroma9 = 9'b000000000;
        12'd84: chroma9 = 9'b000000000;
        12'd85: chroma9 = 9'b000000000;
        12'd86: chroma9 = 9'b000000000;
        12'd87: chroma9 = 9'b000000000;
        12'd88: chroma9 = 9'b000000000;
        12'd89: chroma9 = 9'b000000000;
        12'd90: chroma9 = 9'b000000000;
        12'd91: chroma9 = 9'b000000000;
        12'd92: chroma9 = 9'b000000000;
        12'd93: chroma9 = 9'b000000000;
        12'd94: chroma9 = 9'b000000000;
        12'd95: chroma9 = 9'b000000000;
        12'd96: chroma9 = 9'b000000000;
        12'd97: chroma9 = 9'b000000000;
        12'd98: chroma9 = 9'b000000000;
        12'd99: chroma9 = 9'b000000000;
        12'd100: chroma9 = 9'b000000000;
        12'd101: chroma9 = 9'b000000000;
        12'd102: chroma9 = 9'b000000000;
        12'd103: chroma9 = 9'b000000000;
        12'd104: chroma9 = 9'b000000000;
        12'd105: chroma9 = 9'b000000000;
        12'd106: chroma9 = 9'b000000000;
        12'd107: chroma9 = 9'b000000000;
        12'd108: chroma9 = 9'b000000000;
        12'd109: chroma9 = 9'b000000000;
        12'd110: chroma9 = 9'b000000000;
        12'd111: chroma9 = 9'b000000000;
        12'd112: chroma9 = 9'b000000000;
        12'd113: chroma9 = 9'b000000000;
        12'd114: chroma9 = 9'b000000000;
        12'd115: chroma9 = 9'b000000000;
        12'd116: chroma9 = 9'b000000000;
        12'd117: chroma9 = 9'b000000000;
        12'd118: chroma9 = 9'b000000000;
        12'd119: chroma9 = 9'b000000000;
        12'd120: chroma9 = 9'b000000000;
        12'd121: chroma9 = 9'b000000000;
        12'd122: chroma9 = 9'b000000000;
        12'd123: chroma9 = 9'b000000000;
        12'd124: chroma9 = 9'b000000000;
        12'd125: chroma9 = 9'b000000000;
        12'd126: chroma9 = 9'b000000000;
        12'd127: chroma9 = 9'b000000000;
        12'd128: chroma9 = 9'b000000000;
        12'd129: chroma9 = 9'b000000000;
        12'd130: chroma9 = 9'b000000000;
        12'd131: chroma9 = 9'b000000000;
        12'd132: chroma9 = 9'b000000000;
        12'd133: chroma9 = 9'b000000000;
        12'd134: chroma9 = 9'b000000000;
        12'd135: chroma9 = 9'b000000000;
        12'd136: chroma9 = 9'b000000000;
        12'd137: chroma9 = 9'b000000000;
        12'd138: chroma9 = 9'b000000000;
        12'd139: chroma9 = 9'b000000000;
        12'd140: chroma9 = 9'b000000000;
        12'd141: chroma9 = 9'b000000000;
        12'd142: chroma9 = 9'b000000000;
        12'd143: chroma9 = 9'b000000000;
        12'd144: chroma9 = 9'b000000000;
        12'd145: chroma9 = 9'b000000000;
        12'd146: chroma9 = 9'b000000000;
        12'd147: chroma9 = 9'b000000000;
        12'd148: chroma9 = 9'b000000000;
        12'd149: chroma9 = 9'b000000000;
        12'd150: chroma9 = 9'b000000000;
        12'd151: chroma9 = 9'b000000000;
        12'd152: chroma9 = 9'b000000000;
        12'd153: chroma9 = 9'b000000000;
        12'd154: chroma9 = 9'b000000000;
        12'd155: chroma9 = 9'b000000000;
        12'd156: chroma9 = 9'b000000000;
        12'd157: chroma9 = 9'b000000000;
        12'd158: chroma9 = 9'b000000000;
        12'd159: chroma9 = 9'b000000000;
        12'd160: chroma9 = 9'b000000000;
        12'd161: chroma9 = 9'b000000000;
        12'd162: chroma9 = 9'b000000000;
        12'd163: chroma9 = 9'b000000000;
        12'd164: chroma9 = 9'b000000000;
        12'd165: chroma9 = 9'b000000000;
        12'd166: chroma9 = 9'b000000000;
        12'd167: chroma9 = 9'b000000000;
        12'd168: chroma9 = 9'b000000000;
        12'd169: chroma9 = 9'b000000000;
        12'd170: chroma9 = 9'b000000000;
        12'd171: chroma9 = 9'b000000000;
        12'd172: chroma9 = 9'b000000000;
        12'd173: chroma9 = 9'b000000000;
        12'd174: chroma9 = 9'b000000000;
        12'd175: chroma9 = 9'b000000000;
        12'd176: chroma9 = 9'b000000000;
        12'd177: chroma9 = 9'b000000000;
        12'd178: chroma9 = 9'b000000000;
        12'd179: chroma9 = 9'b000000000;
        12'd180: chroma9 = 9'b000000000;
        12'd181: chroma9 = 9'b000000000;
        12'd182: chroma9 = 9'b000000000;
        12'd183: chroma9 = 9'b000000000;
        12'd184: chroma9 = 9'b000000000;
        12'd185: chroma9 = 9'b000000000;
        12'd186: chroma9 = 9'b000000000;
        12'd187: chroma9 = 9'b000000000;
        12'd188: chroma9 = 9'b000000000;
        12'd189: chroma9 = 9'b000000000;
        12'd190: chroma9 = 9'b000000000;
        12'd191: chroma9 = 9'b000000000;
        12'd192: chroma9 = 9'b000000000;
        12'd193: chroma9 = 9'b000000000;
        12'd194: chroma9 = 9'b000000000;
        12'd195: chroma9 = 9'b000000000;
        12'd196: chroma9 = 9'b000000000;
        12'd197: chroma9 = 9'b000000000;
        12'd198: chroma9 = 9'b000000000;
        12'd199: chroma9 = 9'b000000000;
        12'd200: chroma9 = 9'b000000000;
        12'd201: chroma9 = 9'b000000000;
        12'd202: chroma9 = 9'b000000000;
        12'd203: chroma9 = 9'b000000000;
        12'd204: chroma9 = 9'b000000000;
        12'd205: chroma9 = 9'b000000000;
        12'd206: chroma9 = 9'b000000000;
        12'd207: chroma9 = 9'b000000000;
        12'd208: chroma9 = 9'b000000000;
        12'd209: chroma9 = 9'b000000000;
        12'd210: chroma9 = 9'b000000000;
        12'd211: chroma9 = 9'b000000000;
        12'd212: chroma9 = 9'b000000000;
        12'd213: chroma9 = 9'b000000000;
        12'd214: chroma9 = 9'b000000000;
        12'd215: chroma9 = 9'b000000000;
        12'd216: chroma9 = 9'b000000000;
        12'd217: chroma9 = 9'b000000000;
        12'd218: chroma9 = 9'b000000000;
        12'd219: chroma9 = 9'b000000000;
        12'd220: chroma9 = 9'b000000000;
        12'd221: chroma9 = 9'b000000000;
        12'd222: chroma9 = 9'b000000000;
        12'd223: chroma9 = 9'b000000000;
        12'd224: chroma9 = 9'b000000000;
        12'd225: chroma9 = 9'b000000000;
        12'd226: chroma9 = 9'b000000000;
        12'd227: chroma9 = 9'b000000000;
        12'd228: chroma9 = 9'b000000000;
        12'd229: chroma9 = 9'b000000000;
        12'd230: chroma9 = 9'b000000000;
        12'd231: chroma9 = 9'b000000000;
        12'd232: chroma9 = 9'b000000000;
        12'd233: chroma9 = 9'b000000000;
        12'd234: chroma9 = 9'b000000000;
        12'd235: chroma9 = 9'b000000000;
        12'd236: chroma9 = 9'b000000000;
        12'd237: chroma9 = 9'b000000000;
        12'd238: chroma9 = 9'b000000000;
        12'd239: chroma9 = 9'b000000000;
        12'd240: chroma9 = 9'b000000000;
        12'd241: chroma9 = 9'b000000000;
        12'd242: chroma9 = 9'b000000000;
        12'd243: chroma9 = 9'b000000000;
        12'd244: chroma9 = 9'b000000000;
        12'd245: chroma9 = 9'b000000000;
        12'd246: chroma9 = 9'b000000000;
        12'd247: chroma9 = 9'b000000000;
        12'd248: chroma9 = 9'b000000000;
        12'd249: chroma9 = 9'b000000000;
        12'd250: chroma9 = 9'b000000000;
        12'd251: chroma9 = 9'b000000000;
        12'd252: chroma9 = 9'b000000000;
        12'd253: chroma9 = 9'b000000000;
        12'd254: chroma9 = 9'b000000000;
        12'd255: chroma9 = 9'b000000000;
        12'd256: chroma9 = 9'b100000000;
        12'd257: chroma9 = 9'b100000000;
        12'd258: chroma9 = 9'b100000001;
        12'd259: chroma9 = 9'b100000010;
        12'd260: chroma9 = 9'b100000011;
        12'd261: chroma9 = 9'b100000100;
        12'd262: chroma9 = 9'b100000101;
        12'd263: chroma9 = 9'b100000110;
        12'd264: chroma9 = 9'b100000111;
        12'd265: chroma9 = 9'b100001000;
        12'd266: chroma9 = 9'b100001001;
        12'd267: chroma9 = 9'b100001010;
        12'd268: chroma9 = 9'b100001011;
        12'd269: chroma9 = 9'b100001100;
        12'd270: chroma9 = 9'b100001101;
        12'd271: chroma9 = 9'b100001110;
        12'd272: chroma9 = 9'b100001111;
        12'd273: chroma9 = 9'b100010000;
        12'd274: chroma9 = 9'b100010001;
        12'd275: chroma9 = 9'b100010001;
        12'd276: chroma9 = 9'b100010010;
        12'd277: chroma9 = 9'b100010011;
        12'd278: chroma9 = 9'b100010100;
        12'd279: chroma9 = 9'b100010101;
        12'd280: chroma9 = 9'b100010110;
        12'd281: chroma9 = 9'b100010111;
        12'd282: chroma9 = 9'b100010111;
        12'd283: chroma9 = 9'b100011000;
        12'd284: chroma9 = 9'b100011001;
        12'd285: chroma9 = 9'b100011010;
        12'd286: chroma9 = 9'b100011010;
        12'd287: chroma9 = 9'b100011011;
        12'd288: chroma9 = 9'b100011100;
        12'd289: chroma9 = 9'b100011100;
        12'd290: chroma9 = 9'b100011101;
        12'd291: chroma9 = 9'b100011110;
        12'd292: chroma9 = 9'b100011110;
        12'd293: chroma9 = 9'b100011111;
        12'd294: chroma9 = 9'b100100000;
        12'd295: chroma9 = 9'b100100000;
        12'd296: chroma9 = 9'b100100001;
        12'd297: chroma9 = 9'b100100001;
        12'd298: chroma9 = 9'b100100010;
        12'd299: chroma9 = 9'b100100010;
        12'd300: chroma9 = 9'b100100011;
        12'd301: chroma9 = 9'b100100011;
        12'd302: chroma9 = 9'b100100100;
        12'd303: chroma9 = 9'b100100100;
        12'd304: chroma9 = 9'b100100100;
        12'd305: chroma9 = 9'b100100101;
        12'd306: chroma9 = 9'b100100101;
        12'd307: chroma9 = 9'b100100101;
        12'd308: chroma9 = 9'b100100110;
        12'd309: chroma9 = 9'b100100110;
        12'd310: chroma9 = 9'b100100110;
        12'd311: chroma9 = 9'b100100111;
        12'd312: chroma9 = 9'b100100111;
        12'd313: chroma9 = 9'b100100111;
        12'd314: chroma9 = 9'b100100111;
        12'd315: chroma9 = 9'b100100111;
        12'd316: chroma9 = 9'b100100111;
        12'd317: chroma9 = 9'b100100111;
        12'd318: chroma9 = 9'b100100111;
        12'd319: chroma9 = 9'b100100111;
        12'd320: chroma9 = 9'b100100111;
        12'd321: chroma9 = 9'b100100111;
        12'd322: chroma9 = 9'b100100111;
        12'd323: chroma9 = 9'b100100111;
        12'd324: chroma9 = 9'b100100111;
        12'd325: chroma9 = 9'b100100111;
        12'd326: chroma9 = 9'b100100111;
        12'd327: chroma9 = 9'b100100111;
        12'd328: chroma9 = 9'b100100111;
        12'd329: chroma9 = 9'b100100111;
        12'd330: chroma9 = 9'b100100110;
        12'd331: chroma9 = 9'b100100110;
        12'd332: chroma9 = 9'b100100110;
        12'd333: chroma9 = 9'b100100101;
        12'd334: chroma9 = 9'b100100101;
        12'd335: chroma9 = 9'b100100101;
        12'd336: chroma9 = 9'b100100100;
        12'd337: chroma9 = 9'b100100100;
        12'd338: chroma9 = 9'b100100100;
        12'd339: chroma9 = 9'b100100011;
        12'd340: chroma9 = 9'b100100011;
        12'd341: chroma9 = 9'b100100010;
        12'd342: chroma9 = 9'b100100010;
        12'd343: chroma9 = 9'b100100001;
        12'd344: chroma9 = 9'b100100001;
        12'd345: chroma9 = 9'b100100000;
        12'd346: chroma9 = 9'b100100000;
        12'd347: chroma9 = 9'b100011111;
        12'd348: chroma9 = 9'b100011110;
        12'd349: chroma9 = 9'b100011110;
        12'd350: chroma9 = 9'b100011101;
        12'd351: chroma9 = 9'b100011100;
        12'd352: chroma9 = 9'b100011100;
        12'd353: chroma9 = 9'b100011011;
        12'd354: chroma9 = 9'b100011010;
        12'd355: chroma9 = 9'b100011010;
        12'd356: chroma9 = 9'b100011001;
        12'd357: chroma9 = 9'b100011000;
        12'd358: chroma9 = 9'b100010111;
        12'd359: chroma9 = 9'b100010111;
        12'd360: chroma9 = 9'b100010110;
        12'd361: chroma9 = 9'b100010101;
        12'd362: chroma9 = 9'b100010100;
        12'd363: chroma9 = 9'b100010011;
        12'd364: chroma9 = 9'b100010010;
        12'd365: chroma9 = 9'b100010001;
        12'd366: chroma9 = 9'b100010001;
        12'd367: chroma9 = 9'b100010000;
        12'd368: chroma9 = 9'b100001111;
        12'd369: chroma9 = 9'b100001110;
        12'd370: chroma9 = 9'b100001101;
        12'd371: chroma9 = 9'b100001100;
        12'd372: chroma9 = 9'b100001011;
        12'd373: chroma9 = 9'b100001010;
        12'd374: chroma9 = 9'b100001001;
        12'd375: chroma9 = 9'b100001000;
        12'd376: chroma9 = 9'b100000111;
        12'd377: chroma9 = 9'b100000110;
        12'd378: chroma9 = 9'b100000101;
        12'd379: chroma9 = 9'b100000100;
        12'd380: chroma9 = 9'b100000011;
        12'd381: chroma9 = 9'b100000010;
        12'd382: chroma9 = 9'b100000001;
        12'd383: chroma9 = 9'b100000000;
        12'd384: chroma9 = 9'b100000000;
        12'd385: chroma9 = 9'b100000000;
        12'd386: chroma9 = 9'b011111111;
        12'd387: chroma9 = 9'b011111110;
        12'd388: chroma9 = 9'b011111101;
        12'd389: chroma9 = 9'b011111100;
        12'd390: chroma9 = 9'b011111011;
        12'd391: chroma9 = 9'b011111010;
        12'd392: chroma9 = 9'b011111001;
        12'd393: chroma9 = 9'b011111000;
        12'd394: chroma9 = 9'b011110111;
        12'd395: chroma9 = 9'b011110110;
        12'd396: chroma9 = 9'b011110101;
        12'd397: chroma9 = 9'b011110100;
        12'd398: chroma9 = 9'b011110011;
        12'd399: chroma9 = 9'b011110010;
        12'd400: chroma9 = 9'b011110001;
        12'd401: chroma9 = 9'b011110000;
        12'd402: chroma9 = 9'b011101111;
        12'd403: chroma9 = 9'b011101111;
        12'd404: chroma9 = 9'b011101110;
        12'd405: chroma9 = 9'b011101101;
        12'd406: chroma9 = 9'b011101100;
        12'd407: chroma9 = 9'b011101011;
        12'd408: chroma9 = 9'b011101010;
        12'd409: chroma9 = 9'b011101001;
        12'd410: chroma9 = 9'b011101001;
        12'd411: chroma9 = 9'b011101000;
        12'd412: chroma9 = 9'b011100111;
        12'd413: chroma9 = 9'b011100110;
        12'd414: chroma9 = 9'b011100110;
        12'd415: chroma9 = 9'b011100101;
        12'd416: chroma9 = 9'b011100100;
        12'd417: chroma9 = 9'b011100100;
        12'd418: chroma9 = 9'b011100011;
        12'd419: chroma9 = 9'b011100010;
        12'd420: chroma9 = 9'b011100010;
        12'd421: chroma9 = 9'b011100001;
        12'd422: chroma9 = 9'b011100000;
        12'd423: chroma9 = 9'b011100000;
        12'd424: chroma9 = 9'b011011111;
        12'd425: chroma9 = 9'b011011111;
        12'd426: chroma9 = 9'b011011110;
        12'd427: chroma9 = 9'b011011110;
        12'd428: chroma9 = 9'b011011101;
        12'd429: chroma9 = 9'b011011101;
        12'd430: chroma9 = 9'b011011100;
        12'd431: chroma9 = 9'b011011100;
        12'd432: chroma9 = 9'b011011100;
        12'd433: chroma9 = 9'b011011011;
        12'd434: chroma9 = 9'b011011011;
        12'd435: chroma9 = 9'b011011011;
        12'd436: chroma9 = 9'b011011010;
        12'd437: chroma9 = 9'b011011010;
        12'd438: chroma9 = 9'b011011010;
        12'd439: chroma9 = 9'b011011001;
        12'd440: chroma9 = 9'b011011001;
        12'd441: chroma9 = 9'b011011001;
        12'd442: chroma9 = 9'b011011001;
        12'd443: chroma9 = 9'b011011001;
        12'd444: chroma9 = 9'b011011001;
        12'd445: chroma9 = 9'b011011001;
        12'd446: chroma9 = 9'b011011001;
        12'd447: chroma9 = 9'b011011001;
        12'd448: chroma9 = 9'b011011001;
        12'd449: chroma9 = 9'b011011001;
        12'd450: chroma9 = 9'b011011001;
        12'd451: chroma9 = 9'b011011001;
        12'd452: chroma9 = 9'b011011001;
        12'd453: chroma9 = 9'b011011001;
        12'd454: chroma9 = 9'b011011001;
        12'd455: chroma9 = 9'b011011001;
        12'd456: chroma9 = 9'b011011001;
        12'd457: chroma9 = 9'b011011001;
        12'd458: chroma9 = 9'b011011010;
        12'd459: chroma9 = 9'b011011010;
        12'd460: chroma9 = 9'b011011010;
        12'd461: chroma9 = 9'b011011011;
        12'd462: chroma9 = 9'b011011011;
        12'd463: chroma9 = 9'b011011011;
        12'd464: chroma9 = 9'b011011100;
        12'd465: chroma9 = 9'b011011100;
        12'd466: chroma9 = 9'b011011100;
        12'd467: chroma9 = 9'b011011101;
        12'd468: chroma9 = 9'b011011101;
        12'd469: chroma9 = 9'b011011110;
        12'd470: chroma9 = 9'b011011110;
        12'd471: chroma9 = 9'b011011111;
        12'd472: chroma9 = 9'b011011111;
        12'd473: chroma9 = 9'b011100000;
        12'd474: chroma9 = 9'b011100000;
        12'd475: chroma9 = 9'b011100001;
        12'd476: chroma9 = 9'b011100010;
        12'd477: chroma9 = 9'b011100010;
        12'd478: chroma9 = 9'b011100011;
        12'd479: chroma9 = 9'b011100100;
        12'd480: chroma9 = 9'b011100100;
        12'd481: chroma9 = 9'b011100101;
        12'd482: chroma9 = 9'b011100110;
        12'd483: chroma9 = 9'b011100110;
        12'd484: chroma9 = 9'b011100111;
        12'd485: chroma9 = 9'b011101000;
        12'd486: chroma9 = 9'b011101001;
        12'd487: chroma9 = 9'b011101001;
        12'd488: chroma9 = 9'b011101010;
        12'd489: chroma9 = 9'b011101011;
        12'd490: chroma9 = 9'b011101100;
        12'd491: chroma9 = 9'b011101101;
        12'd492: chroma9 = 9'b011101110;
        12'd493: chroma9 = 9'b011101111;
        12'd494: chroma9 = 9'b011101111;
        12'd495: chroma9 = 9'b011110000;
        12'd496: chroma9 = 9'b011110001;
        12'd497: chroma9 = 9'b011110010;
        12'd498: chroma9 = 9'b011110011;
        12'd499: chroma9 = 9'b011110100;
        12'd500: chroma9 = 9'b011110101;
        12'd501: chroma9 = 9'b011110110;
        12'd502: chroma9 = 9'b011110111;
        12'd503: chroma9 = 9'b011111000;
        12'd504: chroma9 = 9'b011111001;
        12'd505: chroma9 = 9'b011111010;
        12'd506: chroma9 = 9'b011111011;
        12'd507: chroma9 = 9'b011111100;
        12'd508: chroma9 = 9'b011111101;
        12'd509: chroma9 = 9'b011111110;
        12'd510: chroma9 = 9'b011111111;
        12'd511: chroma9 = 9'b100000000;
        12'd512: chroma9 = 9'b100000000;
        12'd513: chroma9 = 9'b100000001;
        12'd514: chroma9 = 9'b100000010;
        12'd515: chroma9 = 9'b100000100;
        12'd516: chroma9 = 9'b100000101;
        12'd517: chroma9 = 9'b100000110;
        12'd518: chroma9 = 9'b100001000;
        12'd519: chroma9 = 9'b100001001;
        12'd520: chroma9 = 9'b100001010;
        12'd521: chroma9 = 9'b100001100;
        12'd522: chroma9 = 9'b100001101;
        12'd523: chroma9 = 9'b100001110;
        12'd524: chroma9 = 9'b100001111;
        12'd525: chroma9 = 9'b100010001;
        12'd526: chroma9 = 9'b100010010;
        12'd527: chroma9 = 9'b100010011;
        12'd528: chroma9 = 9'b100010101;
        12'd529: chroma9 = 9'b100010110;
        12'd530: chroma9 = 9'b100010111;
        12'd531: chroma9 = 9'b100011000;
        12'd532: chroma9 = 9'b100011001;
        12'd533: chroma9 = 9'b100011011;
        12'd534: chroma9 = 9'b100011100;
        12'd535: chroma9 = 9'b100011101;
        12'd536: chroma9 = 9'b100011110;
        12'd537: chroma9 = 9'b100011111;
        12'd538: chroma9 = 9'b100100000;
        12'd539: chroma9 = 9'b100100001;
        12'd540: chroma9 = 9'b100100010;
        12'd541: chroma9 = 9'b100100011;
        12'd542: chroma9 = 9'b100100100;
        12'd543: chroma9 = 9'b100100101;
        12'd544: chroma9 = 9'b100100110;
        12'd545: chroma9 = 9'b100100111;
        12'd546: chroma9 = 9'b100101000;
        12'd547: chroma9 = 9'b100101001;
        12'd548: chroma9 = 9'b100101010;
        12'd549: chroma9 = 9'b100101011;
        12'd550: chroma9 = 9'b100101100;
        12'd551: chroma9 = 9'b100101100;
        12'd552: chroma9 = 9'b100101101;
        12'd553: chroma9 = 9'b100101110;
        12'd554: chroma9 = 9'b100101111;
        12'd555: chroma9 = 9'b100101111;
        12'd556: chroma9 = 9'b100110000;
        12'd557: chroma9 = 9'b100110001;
        12'd558: chroma9 = 9'b100110001;
        12'd559: chroma9 = 9'b100110010;
        12'd560: chroma9 = 9'b100110010;
        12'd561: chroma9 = 9'b100110011;
        12'd562: chroma9 = 9'b100110011;
        12'd563: chroma9 = 9'b100110100;
        12'd564: chroma9 = 9'b100110100;
        12'd565: chroma9 = 9'b100110101;
        12'd566: chroma9 = 9'b100110101;
        12'd567: chroma9 = 9'b100110101;
        12'd568: chroma9 = 9'b100110101;
        12'd569: chroma9 = 9'b100110110;
        12'd570: chroma9 = 9'b100110110;
        12'd571: chroma9 = 9'b100110110;
        12'd572: chroma9 = 9'b100110110;
        12'd573: chroma9 = 9'b100110110;
        12'd574: chroma9 = 9'b100110110;
        12'd575: chroma9 = 9'b100110110;
        12'd576: chroma9 = 9'b100110110;
        12'd577: chroma9 = 9'b100110110;
        12'd578: chroma9 = 9'b100110110;
        12'd579: chroma9 = 9'b100110110;
        12'd580: chroma9 = 9'b100110110;
        12'd581: chroma9 = 9'b100110110;
        12'd582: chroma9 = 9'b100110110;
        12'd583: chroma9 = 9'b100110110;
        12'd584: chroma9 = 9'b100110101;
        12'd585: chroma9 = 9'b100110101;
        12'd586: chroma9 = 9'b100110101;
        12'd587: chroma9 = 9'b100110101;
        12'd588: chroma9 = 9'b100110100;
        12'd589: chroma9 = 9'b100110100;
        12'd590: chroma9 = 9'b100110011;
        12'd591: chroma9 = 9'b100110011;
        12'd592: chroma9 = 9'b100110010;
        12'd593: chroma9 = 9'b100110010;
        12'd594: chroma9 = 9'b100110001;
        12'd595: chroma9 = 9'b100110001;
        12'd596: chroma9 = 9'b100110000;
        12'd597: chroma9 = 9'b100101111;
        12'd598: chroma9 = 9'b100101111;
        12'd599: chroma9 = 9'b100101110;
        12'd600: chroma9 = 9'b100101101;
        12'd601: chroma9 = 9'b100101100;
        12'd602: chroma9 = 9'b100101100;
        12'd603: chroma9 = 9'b100101011;
        12'd604: chroma9 = 9'b100101010;
        12'd605: chroma9 = 9'b100101001;
        12'd606: chroma9 = 9'b100101000;
        12'd607: chroma9 = 9'b100100111;
        12'd608: chroma9 = 9'b100100110;
        12'd609: chroma9 = 9'b100100101;
        12'd610: chroma9 = 9'b100100100;
        12'd611: chroma9 = 9'b100100011;
        12'd612: chroma9 = 9'b100100010;
        12'd613: chroma9 = 9'b100100001;
        12'd614: chroma9 = 9'b100100000;
        12'd615: chroma9 = 9'b100011111;
        12'd616: chroma9 = 9'b100011110;
        12'd617: chroma9 = 9'b100011101;
        12'd618: chroma9 = 9'b100011100;
        12'd619: chroma9 = 9'b100011011;
        12'd620: chroma9 = 9'b100011001;
        12'd621: chroma9 = 9'b100011000;
        12'd622: chroma9 = 9'b100010111;
        12'd623: chroma9 = 9'b100010110;
        12'd624: chroma9 = 9'b100010101;
        12'd625: chroma9 = 9'b100010011;
        12'd626: chroma9 = 9'b100010010;
        12'd627: chroma9 = 9'b100010001;
        12'd628: chroma9 = 9'b100001111;
        12'd629: chroma9 = 9'b100001110;
        12'd630: chroma9 = 9'b100001101;
        12'd631: chroma9 = 9'b100001100;
        12'd632: chroma9 = 9'b100001010;
        12'd633: chroma9 = 9'b100001001;
        12'd634: chroma9 = 9'b100001000;
        12'd635: chroma9 = 9'b100000110;
        12'd636: chroma9 = 9'b100000101;
        12'd637: chroma9 = 9'b100000100;
        12'd638: chroma9 = 9'b100000010;
        12'd639: chroma9 = 9'b100000001;
        12'd640: chroma9 = 9'b100000000;
        12'd641: chroma9 = 9'b011111111;
        12'd642: chroma9 = 9'b011111110;
        12'd643: chroma9 = 9'b011111100;
        12'd644: chroma9 = 9'b011111011;
        12'd645: chroma9 = 9'b011111010;
        12'd646: chroma9 = 9'b011111000;
        12'd647: chroma9 = 9'b011110111;
        12'd648: chroma9 = 9'b011110110;
        12'd649: chroma9 = 9'b011110100;
        12'd650: chroma9 = 9'b011110011;
        12'd651: chroma9 = 9'b011110010;
        12'd652: chroma9 = 9'b011110001;
        12'd653: chroma9 = 9'b011101111;
        12'd654: chroma9 = 9'b011101110;
        12'd655: chroma9 = 9'b011101101;
        12'd656: chroma9 = 9'b011101011;
        12'd657: chroma9 = 9'b011101010;
        12'd658: chroma9 = 9'b011101001;
        12'd659: chroma9 = 9'b011101000;
        12'd660: chroma9 = 9'b011100111;
        12'd661: chroma9 = 9'b011100101;
        12'd662: chroma9 = 9'b011100100;
        12'd663: chroma9 = 9'b011100011;
        12'd664: chroma9 = 9'b011100010;
        12'd665: chroma9 = 9'b011100001;
        12'd666: chroma9 = 9'b011100000;
        12'd667: chroma9 = 9'b011011111;
        12'd668: chroma9 = 9'b011011110;
        12'd669: chroma9 = 9'b011011101;
        12'd670: chroma9 = 9'b011011100;
        12'd671: chroma9 = 9'b011011011;
        12'd672: chroma9 = 9'b011011010;
        12'd673: chroma9 = 9'b011011001;
        12'd674: chroma9 = 9'b011011000;
        12'd675: chroma9 = 9'b011010111;
        12'd676: chroma9 = 9'b011010110;
        12'd677: chroma9 = 9'b011010101;
        12'd678: chroma9 = 9'b011010100;
        12'd679: chroma9 = 9'b011010100;
        12'd680: chroma9 = 9'b011010011;
        12'd681: chroma9 = 9'b011010010;
        12'd682: chroma9 = 9'b011010001;
        12'd683: chroma9 = 9'b011010001;
        12'd684: chroma9 = 9'b011010000;
        12'd685: chroma9 = 9'b011001111;
        12'd686: chroma9 = 9'b011001111;
        12'd687: chroma9 = 9'b011001110;
        12'd688: chroma9 = 9'b011001110;
        12'd689: chroma9 = 9'b011001101;
        12'd690: chroma9 = 9'b011001101;
        12'd691: chroma9 = 9'b011001100;
        12'd692: chroma9 = 9'b011001100;
        12'd693: chroma9 = 9'b011001011;
        12'd694: chroma9 = 9'b011001011;
        12'd695: chroma9 = 9'b011001011;
        12'd696: chroma9 = 9'b011001011;
        12'd697: chroma9 = 9'b011001010;
        12'd698: chroma9 = 9'b011001010;
        12'd699: chroma9 = 9'b011001010;
        12'd700: chroma9 = 9'b011001010;
        12'd701: chroma9 = 9'b011001010;
        12'd702: chroma9 = 9'b011001010;
        12'd703: chroma9 = 9'b011001010;
        12'd704: chroma9 = 9'b011001010;
        12'd705: chroma9 = 9'b011001010;
        12'd706: chroma9 = 9'b011001010;
        12'd707: chroma9 = 9'b011001010;
        12'd708: chroma9 = 9'b011001010;
        12'd709: chroma9 = 9'b011001010;
        12'd710: chroma9 = 9'b011001010;
        12'd711: chroma9 = 9'b011001010;
        12'd712: chroma9 = 9'b011001011;
        12'd713: chroma9 = 9'b011001011;
        12'd714: chroma9 = 9'b011001011;
        12'd715: chroma9 = 9'b011001011;
        12'd716: chroma9 = 9'b011001100;
        12'd717: chroma9 = 9'b011001100;
        12'd718: chroma9 = 9'b011001101;
        12'd719: chroma9 = 9'b011001101;
        12'd720: chroma9 = 9'b011001110;
        12'd721: chroma9 = 9'b011001110;
        12'd722: chroma9 = 9'b011001111;
        12'd723: chroma9 = 9'b011001111;
        12'd724: chroma9 = 9'b011010000;
        12'd725: chroma9 = 9'b011010001;
        12'd726: chroma9 = 9'b011010001;
        12'd727: chroma9 = 9'b011010010;
        12'd728: chroma9 = 9'b011010011;
        12'd729: chroma9 = 9'b011010100;
        12'd730: chroma9 = 9'b011010100;
        12'd731: chroma9 = 9'b011010101;
        12'd732: chroma9 = 9'b011010110;
        12'd733: chroma9 = 9'b011010111;
        12'd734: chroma9 = 9'b011011000;
        12'd735: chroma9 = 9'b011011001;
        12'd736: chroma9 = 9'b011011010;
        12'd737: chroma9 = 9'b011011011;
        12'd738: chroma9 = 9'b011011100;
        12'd739: chroma9 = 9'b011011101;
        12'd740: chroma9 = 9'b011011110;
        12'd741: chroma9 = 9'b011011111;
        12'd742: chroma9 = 9'b011100000;
        12'd743: chroma9 = 9'b011100001;
        12'd744: chroma9 = 9'b011100010;
        12'd745: chroma9 = 9'b011100011;
        12'd746: chroma9 = 9'b011100100;
        12'd747: chroma9 = 9'b011100101;
        12'd748: chroma9 = 9'b011100111;
        12'd749: chroma9 = 9'b011101000;
        12'd750: chroma9 = 9'b011101001;
        12'd751: chroma9 = 9'b011101010;
        12'd752: chroma9 = 9'b011101011;
        12'd753: chroma9 = 9'b011101101;
        12'd754: chroma9 = 9'b011101110;
        12'd755: chroma9 = 9'b011101111;
        12'd756: chroma9 = 9'b011110001;
        12'd757: chroma9 = 9'b011110010;
        12'd758: chroma9 = 9'b011110011;
        12'd759: chroma9 = 9'b011110100;
        12'd760: chroma9 = 9'b011110110;
        12'd761: chroma9 = 9'b011110111;
        12'd762: chroma9 = 9'b011111000;
        12'd763: chroma9 = 9'b011111010;
        12'd764: chroma9 = 9'b011111011;
        12'd765: chroma9 = 9'b011111100;
        12'd766: chroma9 = 9'b011111110;
        12'd767: chroma9 = 9'b011111111;
        12'd768: chroma9 = 9'b100000000;
        12'd769: chroma9 = 9'b100000001;
        12'd770: chroma9 = 9'b100000011;
        12'd771: chroma9 = 9'b100000101;
        12'd772: chroma9 = 9'b100000110;
        12'd773: chroma9 = 9'b100001000;
        12'd774: chroma9 = 9'b100001010;
        12'd775: chroma9 = 9'b100001011;
        12'd776: chroma9 = 9'b100001101;
        12'd777: chroma9 = 9'b100001111;
        12'd778: chroma9 = 9'b100010001;
        12'd779: chroma9 = 9'b100010010;
        12'd780: chroma9 = 9'b100010100;
        12'd781: chroma9 = 9'b100010101;
        12'd782: chroma9 = 9'b100010111;
        12'd783: chroma9 = 9'b100011001;
        12'd784: chroma9 = 9'b100011010;
        12'd785: chroma9 = 9'b100011100;
        12'd786: chroma9 = 9'b100011101;
        12'd787: chroma9 = 9'b100011111;
        12'd788: chroma9 = 9'b100100000;
        12'd789: chroma9 = 9'b100100010;
        12'd790: chroma9 = 9'b100100011;
        12'd791: chroma9 = 9'b100100101;
        12'd792: chroma9 = 9'b100100110;
        12'd793: chroma9 = 9'b100101000;
        12'd794: chroma9 = 9'b100101001;
        12'd795: chroma9 = 9'b100101011;
        12'd796: chroma9 = 9'b100101100;
        12'd797: chroma9 = 9'b100101101;
        12'd798: chroma9 = 9'b100101111;
        12'd799: chroma9 = 9'b100110000;
        12'd800: chroma9 = 9'b100110001;
        12'd801: chroma9 = 9'b100110010;
        12'd802: chroma9 = 9'b100110011;
        12'd803: chroma9 = 9'b100110101;
        12'd804: chroma9 = 9'b100110110;
        12'd805: chroma9 = 9'b100110111;
        12'd806: chroma9 = 9'b100111000;
        12'd807: chroma9 = 9'b100111001;
        12'd808: chroma9 = 9'b100111010;
        12'd809: chroma9 = 9'b100111011;
        12'd810: chroma9 = 9'b100111100;
        12'd811: chroma9 = 9'b100111100;
        12'd812: chroma9 = 9'b100111101;
        12'd813: chroma9 = 9'b100111110;
        12'd814: chroma9 = 9'b100111111;
        12'd815: chroma9 = 9'b100111111;
        12'd816: chroma9 = 9'b101000000;
        12'd817: chroma9 = 9'b101000001;
        12'd818: chroma9 = 9'b101000001;
        12'd819: chroma9 = 9'b101000010;
        12'd820: chroma9 = 9'b101000010;
        12'd821: chroma9 = 9'b101000011;
        12'd822: chroma9 = 9'b101000011;
        12'd823: chroma9 = 9'b101000100;
        12'd824: chroma9 = 9'b101000100;
        12'd825: chroma9 = 9'b101000100;
        12'd826: chroma9 = 9'b101000101;
        12'd827: chroma9 = 9'b101000101;
        12'd828: chroma9 = 9'b101000101;
        12'd829: chroma9 = 9'b101000101;
        12'd830: chroma9 = 9'b101000101;
        12'd831: chroma9 = 9'b101000101;
        12'd832: chroma9 = 9'b101000101;
        12'd833: chroma9 = 9'b101000101;
        12'd834: chroma9 = 9'b101000101;
        12'd835: chroma9 = 9'b101000101;
        12'd836: chroma9 = 9'b101000101;
        12'd837: chroma9 = 9'b101000101;
        12'd838: chroma9 = 9'b101000101;
        12'd839: chroma9 = 9'b101000100;
        12'd840: chroma9 = 9'b101000100;
        12'd841: chroma9 = 9'b101000100;
        12'd842: chroma9 = 9'b101000011;
        12'd843: chroma9 = 9'b101000011;
        12'd844: chroma9 = 9'b101000010;
        12'd845: chroma9 = 9'b101000010;
        12'd846: chroma9 = 9'b101000001;
        12'd847: chroma9 = 9'b101000001;
        12'd848: chroma9 = 9'b101000000;
        12'd849: chroma9 = 9'b100111111;
        12'd850: chroma9 = 9'b100111111;
        12'd851: chroma9 = 9'b100111110;
        12'd852: chroma9 = 9'b100111101;
        12'd853: chroma9 = 9'b100111100;
        12'd854: chroma9 = 9'b100111100;
        12'd855: chroma9 = 9'b100111011;
        12'd856: chroma9 = 9'b100111010;
        12'd857: chroma9 = 9'b100111001;
        12'd858: chroma9 = 9'b100111000;
        12'd859: chroma9 = 9'b100110111;
        12'd860: chroma9 = 9'b100110110;
        12'd861: chroma9 = 9'b100110101;
        12'd862: chroma9 = 9'b100110011;
        12'd863: chroma9 = 9'b100110010;
        12'd864: chroma9 = 9'b100110001;
        12'd865: chroma9 = 9'b100110000;
        12'd866: chroma9 = 9'b100101111;
        12'd867: chroma9 = 9'b100101101;
        12'd868: chroma9 = 9'b100101100;
        12'd869: chroma9 = 9'b100101011;
        12'd870: chroma9 = 9'b100101001;
        12'd871: chroma9 = 9'b100101000;
        12'd872: chroma9 = 9'b100100110;
        12'd873: chroma9 = 9'b100100101;
        12'd874: chroma9 = 9'b100100011;
        12'd875: chroma9 = 9'b100100010;
        12'd876: chroma9 = 9'b100100000;
        12'd877: chroma9 = 9'b100011111;
        12'd878: chroma9 = 9'b100011101;
        12'd879: chroma9 = 9'b100011100;
        12'd880: chroma9 = 9'b100011010;
        12'd881: chroma9 = 9'b100011001;
        12'd882: chroma9 = 9'b100010111;
        12'd883: chroma9 = 9'b100010101;
        12'd884: chroma9 = 9'b100010100;
        12'd885: chroma9 = 9'b100010010;
        12'd886: chroma9 = 9'b100010001;
        12'd887: chroma9 = 9'b100001111;
        12'd888: chroma9 = 9'b100001101;
        12'd889: chroma9 = 9'b100001011;
        12'd890: chroma9 = 9'b100001010;
        12'd891: chroma9 = 9'b100001000;
        12'd892: chroma9 = 9'b100000110;
        12'd893: chroma9 = 9'b100000101;
        12'd894: chroma9 = 9'b100000011;
        12'd895: chroma9 = 9'b100000001;
        12'd896: chroma9 = 9'b100000000;
        12'd897: chroma9 = 9'b011111111;
        12'd898: chroma9 = 9'b011111101;
        12'd899: chroma9 = 9'b011111011;
        12'd900: chroma9 = 9'b011111010;
        12'd901: chroma9 = 9'b011111000;
        12'd902: chroma9 = 9'b011110110;
        12'd903: chroma9 = 9'b011110101;
        12'd904: chroma9 = 9'b011110011;
        12'd905: chroma9 = 9'b011110001;
        12'd906: chroma9 = 9'b011101111;
        12'd907: chroma9 = 9'b011101110;
        12'd908: chroma9 = 9'b011101100;
        12'd909: chroma9 = 9'b011101011;
        12'd910: chroma9 = 9'b011101001;
        12'd911: chroma9 = 9'b011100111;
        12'd912: chroma9 = 9'b011100110;
        12'd913: chroma9 = 9'b011100100;
        12'd914: chroma9 = 9'b011100011;
        12'd915: chroma9 = 9'b011100001;
        12'd916: chroma9 = 9'b011100000;
        12'd917: chroma9 = 9'b011011110;
        12'd918: chroma9 = 9'b011011101;
        12'd919: chroma9 = 9'b011011011;
        12'd920: chroma9 = 9'b011011010;
        12'd921: chroma9 = 9'b011011000;
        12'd922: chroma9 = 9'b011010111;
        12'd923: chroma9 = 9'b011010101;
        12'd924: chroma9 = 9'b011010100;
        12'd925: chroma9 = 9'b011010011;
        12'd926: chroma9 = 9'b011010001;
        12'd927: chroma9 = 9'b011010000;
        12'd928: chroma9 = 9'b011001111;
        12'd929: chroma9 = 9'b011001110;
        12'd930: chroma9 = 9'b011001101;
        12'd931: chroma9 = 9'b011001011;
        12'd932: chroma9 = 9'b011001010;
        12'd933: chroma9 = 9'b011001001;
        12'd934: chroma9 = 9'b011001000;
        12'd935: chroma9 = 9'b011000111;
        12'd936: chroma9 = 9'b011000110;
        12'd937: chroma9 = 9'b011000101;
        12'd938: chroma9 = 9'b011000100;
        12'd939: chroma9 = 9'b011000100;
        12'd940: chroma9 = 9'b011000011;
        12'd941: chroma9 = 9'b011000010;
        12'd942: chroma9 = 9'b011000001;
        12'd943: chroma9 = 9'b011000001;
        12'd944: chroma9 = 9'b011000000;
        12'd945: chroma9 = 9'b010111111;
        12'd946: chroma9 = 9'b010111111;
        12'd947: chroma9 = 9'b010111110;
        12'd948: chroma9 = 9'b010111110;
        12'd949: chroma9 = 9'b010111101;
        12'd950: chroma9 = 9'b010111101;
        12'd951: chroma9 = 9'b010111100;
        12'd952: chroma9 = 9'b010111100;
        12'd953: chroma9 = 9'b010111100;
        12'd954: chroma9 = 9'b010111011;
        12'd955: chroma9 = 9'b010111011;
        12'd956: chroma9 = 9'b010111011;
        12'd957: chroma9 = 9'b010111011;
        12'd958: chroma9 = 9'b010111011;
        12'd959: chroma9 = 9'b010111011;
        12'd960: chroma9 = 9'b010111011;
        12'd961: chroma9 = 9'b010111011;
        12'd962: chroma9 = 9'b010111011;
        12'd963: chroma9 = 9'b010111011;
        12'd964: chroma9 = 9'b010111011;
        12'd965: chroma9 = 9'b010111011;
        12'd966: chroma9 = 9'b010111011;
        12'd967: chroma9 = 9'b010111100;
        12'd968: chroma9 = 9'b010111100;
        12'd969: chroma9 = 9'b010111100;
        12'd970: chroma9 = 9'b010111101;
        12'd971: chroma9 = 9'b010111101;
        12'd972: chroma9 = 9'b010111110;
        12'd973: chroma9 = 9'b010111110;
        12'd974: chroma9 = 9'b010111111;
        12'd975: chroma9 = 9'b010111111;
        12'd976: chroma9 = 9'b011000000;
        12'd977: chroma9 = 9'b011000001;
        12'd978: chroma9 = 9'b011000001;
        12'd979: chroma9 = 9'b011000010;
        12'd980: chroma9 = 9'b011000011;
        12'd981: chroma9 = 9'b011000100;
        12'd982: chroma9 = 9'b011000100;
        12'd983: chroma9 = 9'b011000101;
        12'd984: chroma9 = 9'b011000110;
        12'd985: chroma9 = 9'b011000111;
        12'd986: chroma9 = 9'b011001000;
        12'd987: chroma9 = 9'b011001001;
        12'd988: chroma9 = 9'b011001010;
        12'd989: chroma9 = 9'b011001011;
        12'd990: chroma9 = 9'b011001101;
        12'd991: chroma9 = 9'b011001110;
        12'd992: chroma9 = 9'b011001111;
        12'd993: chroma9 = 9'b011010000;
        12'd994: chroma9 = 9'b011010001;
        12'd995: chroma9 = 9'b011010011;
        12'd996: chroma9 = 9'b011010100;
        12'd997: chroma9 = 9'b011010101;
        12'd998: chroma9 = 9'b011010111;
        12'd999: chroma9 = 9'b011011000;
        12'd1000: chroma9 = 9'b011011010;
        12'd1001: chroma9 = 9'b011011011;
        12'd1002: chroma9 = 9'b011011101;
        12'd1003: chroma9 = 9'b011011110;
        12'd1004: chroma9 = 9'b011100000;
        12'd1005: chroma9 = 9'b011100001;
        12'd1006: chroma9 = 9'b011100011;
        12'd1007: chroma9 = 9'b011100100;
        12'd1008: chroma9 = 9'b011100110;
        12'd1009: chroma9 = 9'b011100111;
        12'd1010: chroma9 = 9'b011101001;
        12'd1011: chroma9 = 9'b011101011;
        12'd1012: chroma9 = 9'b011101100;
        12'd1013: chroma9 = 9'b011101110;
        12'd1014: chroma9 = 9'b011101111;
        12'd1015: chroma9 = 9'b011110001;
        12'd1016: chroma9 = 9'b011110011;
        12'd1017: chroma9 = 9'b011110101;
        12'd1018: chroma9 = 9'b011110110;
        12'd1019: chroma9 = 9'b011111000;
        12'd1020: chroma9 = 9'b011111010;
        12'd1021: chroma9 = 9'b011111011;
        12'd1022: chroma9 = 9'b011111101;
        12'd1023: chroma9 = 9'b011111111;
        12'd1024: chroma9 = 9'b100000000;
        12'd1025: chroma9 = 9'b100000010;
        12'd1026: chroma9 = 9'b100000100;
        12'd1027: chroma9 = 9'b100000110;
        12'd1028: chroma9 = 9'b100001000;
        12'd1029: chroma9 = 9'b100001010;
        12'd1030: chroma9 = 9'b100001100;
        12'd1031: chroma9 = 9'b100001110;
        12'd1032: chroma9 = 9'b100010000;
        12'd1033: chroma9 = 9'b100010010;
        12'd1034: chroma9 = 9'b100010100;
        12'd1035: chroma9 = 9'b100010110;
        12'd1036: chroma9 = 9'b100011000;
        12'd1037: chroma9 = 9'b100011010;
        12'd1038: chroma9 = 9'b100011100;
        12'd1039: chroma9 = 9'b100011110;
        12'd1040: chroma9 = 9'b100100000;
        12'd1041: chroma9 = 9'b100100010;
        12'd1042: chroma9 = 9'b100100100;
        12'd1043: chroma9 = 9'b100100110;
        12'd1044: chroma9 = 9'b100101000;
        12'd1045: chroma9 = 9'b100101001;
        12'd1046: chroma9 = 9'b100101011;
        12'd1047: chroma9 = 9'b100101101;
        12'd1048: chroma9 = 9'b100101111;
        12'd1049: chroma9 = 9'b100110000;
        12'd1050: chroma9 = 9'b100110010;
        12'd1051: chroma9 = 9'b100110100;
        12'd1052: chroma9 = 9'b100110101;
        12'd1053: chroma9 = 9'b100110111;
        12'd1054: chroma9 = 9'b100111001;
        12'd1055: chroma9 = 9'b100111010;
        12'd1056: chroma9 = 9'b100111100;
        12'd1057: chroma9 = 9'b100111101;
        12'd1058: chroma9 = 9'b100111110;
        12'd1059: chroma9 = 9'b101000000;
        12'd1060: chroma9 = 9'b101000001;
        12'd1061: chroma9 = 9'b101000011;
        12'd1062: chroma9 = 9'b101000100;
        12'd1063: chroma9 = 9'b101000101;
        12'd1064: chroma9 = 9'b101000110;
        12'd1065: chroma9 = 9'b101000111;
        12'd1066: chroma9 = 9'b101001000;
        12'd1067: chroma9 = 9'b101001001;
        12'd1068: chroma9 = 9'b101001010;
        12'd1069: chroma9 = 9'b101001011;
        12'd1070: chroma9 = 9'b101001100;
        12'd1071: chroma9 = 9'b101001101;
        12'd1072: chroma9 = 9'b101001110;
        12'd1073: chroma9 = 9'b101001111;
        12'd1074: chroma9 = 9'b101010000;
        12'd1075: chroma9 = 9'b101010000;
        12'd1076: chroma9 = 9'b101010001;
        12'd1077: chroma9 = 9'b101010001;
        12'd1078: chroma9 = 9'b101010010;
        12'd1079: chroma9 = 9'b101010010;
        12'd1080: chroma9 = 9'b101010011;
        12'd1081: chroma9 = 9'b101010011;
        12'd1082: chroma9 = 9'b101010100;
        12'd1083: chroma9 = 9'b101010100;
        12'd1084: chroma9 = 9'b101010100;
        12'd1085: chroma9 = 9'b101010100;
        12'd1086: chroma9 = 9'b101010100;
        12'd1087: chroma9 = 9'b101010100;
        12'd1088: chroma9 = 9'b101010100;
        12'd1089: chroma9 = 9'b101010100;
        12'd1090: chroma9 = 9'b101010100;
        12'd1091: chroma9 = 9'b101010100;
        12'd1092: chroma9 = 9'b101010100;
        12'd1093: chroma9 = 9'b101010100;
        12'd1094: chroma9 = 9'b101010100;
        12'd1095: chroma9 = 9'b101010011;
        12'd1096: chroma9 = 9'b101010011;
        12'd1097: chroma9 = 9'b101010010;
        12'd1098: chroma9 = 9'b101010010;
        12'd1099: chroma9 = 9'b101010001;
        12'd1100: chroma9 = 9'b101010001;
        12'd1101: chroma9 = 9'b101010000;
        12'd1102: chroma9 = 9'b101010000;
        12'd1103: chroma9 = 9'b101001111;
        12'd1104: chroma9 = 9'b101001110;
        12'd1105: chroma9 = 9'b101001101;
        12'd1106: chroma9 = 9'b101001100;
        12'd1107: chroma9 = 9'b101001011;
        12'd1108: chroma9 = 9'b101001010;
        12'd1109: chroma9 = 9'b101001001;
        12'd1110: chroma9 = 9'b101001000;
        12'd1111: chroma9 = 9'b101000111;
        12'd1112: chroma9 = 9'b101000110;
        12'd1113: chroma9 = 9'b101000101;
        12'd1114: chroma9 = 9'b101000100;
        12'd1115: chroma9 = 9'b101000011;
        12'd1116: chroma9 = 9'b101000001;
        12'd1117: chroma9 = 9'b101000000;
        12'd1118: chroma9 = 9'b100111110;
        12'd1119: chroma9 = 9'b100111101;
        12'd1120: chroma9 = 9'b100111100;
        12'd1121: chroma9 = 9'b100111010;
        12'd1122: chroma9 = 9'b100111001;
        12'd1123: chroma9 = 9'b100110111;
        12'd1124: chroma9 = 9'b100110101;
        12'd1125: chroma9 = 9'b100110100;
        12'd1126: chroma9 = 9'b100110010;
        12'd1127: chroma9 = 9'b100110000;
        12'd1128: chroma9 = 9'b100101111;
        12'd1129: chroma9 = 9'b100101101;
        12'd1130: chroma9 = 9'b100101011;
        12'd1131: chroma9 = 9'b100101001;
        12'd1132: chroma9 = 9'b100101000;
        12'd1133: chroma9 = 9'b100100110;
        12'd1134: chroma9 = 9'b100100100;
        12'd1135: chroma9 = 9'b100100010;
        12'd1136: chroma9 = 9'b100100000;
        12'd1137: chroma9 = 9'b100011110;
        12'd1138: chroma9 = 9'b100011100;
        12'd1139: chroma9 = 9'b100011010;
        12'd1140: chroma9 = 9'b100011000;
        12'd1141: chroma9 = 9'b100010110;
        12'd1142: chroma9 = 9'b100010100;
        12'd1143: chroma9 = 9'b100010010;
        12'd1144: chroma9 = 9'b100010000;
        12'd1145: chroma9 = 9'b100001110;
        12'd1146: chroma9 = 9'b100001100;
        12'd1147: chroma9 = 9'b100001010;
        12'd1148: chroma9 = 9'b100001000;
        12'd1149: chroma9 = 9'b100000110;
        12'd1150: chroma9 = 9'b100000100;
        12'd1151: chroma9 = 9'b100000010;
        12'd1152: chroma9 = 9'b100000000;
        12'd1153: chroma9 = 9'b011111110;
        12'd1154: chroma9 = 9'b011111100;
        12'd1155: chroma9 = 9'b011111010;
        12'd1156: chroma9 = 9'b011111000;
        12'd1157: chroma9 = 9'b011110110;
        12'd1158: chroma9 = 9'b011110100;
        12'd1159: chroma9 = 9'b011110010;
        12'd1160: chroma9 = 9'b011110000;
        12'd1161: chroma9 = 9'b011101110;
        12'd1162: chroma9 = 9'b011101100;
        12'd1163: chroma9 = 9'b011101010;
        12'd1164: chroma9 = 9'b011101000;
        12'd1165: chroma9 = 9'b011100110;
        12'd1166: chroma9 = 9'b011100100;
        12'd1167: chroma9 = 9'b011100010;
        12'd1168: chroma9 = 9'b011100000;
        12'd1169: chroma9 = 9'b011011110;
        12'd1170: chroma9 = 9'b011011100;
        12'd1171: chroma9 = 9'b011011010;
        12'd1172: chroma9 = 9'b011011000;
        12'd1173: chroma9 = 9'b011010111;
        12'd1174: chroma9 = 9'b011010101;
        12'd1175: chroma9 = 9'b011010011;
        12'd1176: chroma9 = 9'b011010001;
        12'd1177: chroma9 = 9'b011010000;
        12'd1178: chroma9 = 9'b011001110;
        12'd1179: chroma9 = 9'b011001100;
        12'd1180: chroma9 = 9'b011001011;
        12'd1181: chroma9 = 9'b011001001;
        12'd1182: chroma9 = 9'b011000111;
        12'd1183: chroma9 = 9'b011000110;
        12'd1184: chroma9 = 9'b011000100;
        12'd1185: chroma9 = 9'b011000011;
        12'd1186: chroma9 = 9'b011000010;
        12'd1187: chroma9 = 9'b011000000;
        12'd1188: chroma9 = 9'b010111111;
        12'd1189: chroma9 = 9'b010111101;
        12'd1190: chroma9 = 9'b010111100;
        12'd1191: chroma9 = 9'b010111011;
        12'd1192: chroma9 = 9'b010111010;
        12'd1193: chroma9 = 9'b010111001;
        12'd1194: chroma9 = 9'b010111000;
        12'd1195: chroma9 = 9'b010110111;
        12'd1196: chroma9 = 9'b010110110;
        12'd1197: chroma9 = 9'b010110101;
        12'd1198: chroma9 = 9'b010110100;
        12'd1199: chroma9 = 9'b010110011;
        12'd1200: chroma9 = 9'b010110010;
        12'd1201: chroma9 = 9'b010110001;
        12'd1202: chroma9 = 9'b010110000;
        12'd1203: chroma9 = 9'b010110000;
        12'd1204: chroma9 = 9'b010101111;
        12'd1205: chroma9 = 9'b010101111;
        12'd1206: chroma9 = 9'b010101110;
        12'd1207: chroma9 = 9'b010101110;
        12'd1208: chroma9 = 9'b010101101;
        12'd1209: chroma9 = 9'b010101101;
        12'd1210: chroma9 = 9'b010101100;
        12'd1211: chroma9 = 9'b010101100;
        12'd1212: chroma9 = 9'b010101100;
        12'd1213: chroma9 = 9'b010101100;
        12'd1214: chroma9 = 9'b010101100;
        12'd1215: chroma9 = 9'b010101100;
        12'd1216: chroma9 = 9'b010101100;
        12'd1217: chroma9 = 9'b010101100;
        12'd1218: chroma9 = 9'b010101100;
        12'd1219: chroma9 = 9'b010101100;
        12'd1220: chroma9 = 9'b010101100;
        12'd1221: chroma9 = 9'b010101100;
        12'd1222: chroma9 = 9'b010101100;
        12'd1223: chroma9 = 9'b010101101;
        12'd1224: chroma9 = 9'b010101101;
        12'd1225: chroma9 = 9'b010101110;
        12'd1226: chroma9 = 9'b010101110;
        12'd1227: chroma9 = 9'b010101111;
        12'd1228: chroma9 = 9'b010101111;
        12'd1229: chroma9 = 9'b010110000;
        12'd1230: chroma9 = 9'b010110000;
        12'd1231: chroma9 = 9'b010110001;
        12'd1232: chroma9 = 9'b010110010;
        12'd1233: chroma9 = 9'b010110011;
        12'd1234: chroma9 = 9'b010110100;
        12'd1235: chroma9 = 9'b010110101;
        12'd1236: chroma9 = 9'b010110110;
        12'd1237: chroma9 = 9'b010110111;
        12'd1238: chroma9 = 9'b010111000;
        12'd1239: chroma9 = 9'b010111001;
        12'd1240: chroma9 = 9'b010111010;
        12'd1241: chroma9 = 9'b010111011;
        12'd1242: chroma9 = 9'b010111100;
        12'd1243: chroma9 = 9'b010111101;
        12'd1244: chroma9 = 9'b010111111;
        12'd1245: chroma9 = 9'b011000000;
        12'd1246: chroma9 = 9'b011000010;
        12'd1247: chroma9 = 9'b011000011;
        12'd1248: chroma9 = 9'b011000100;
        12'd1249: chroma9 = 9'b011000110;
        12'd1250: chroma9 = 9'b011000111;
        12'd1251: chroma9 = 9'b011001001;
        12'd1252: chroma9 = 9'b011001011;
        12'd1253: chroma9 = 9'b011001100;
        12'd1254: chroma9 = 9'b011001110;
        12'd1255: chroma9 = 9'b011010000;
        12'd1256: chroma9 = 9'b011010001;
        12'd1257: chroma9 = 9'b011010011;
        12'd1258: chroma9 = 9'b011010101;
        12'd1259: chroma9 = 9'b011010111;
        12'd1260: chroma9 = 9'b011011000;
        12'd1261: chroma9 = 9'b011011010;
        12'd1262: chroma9 = 9'b011011100;
        12'd1263: chroma9 = 9'b011011110;
        12'd1264: chroma9 = 9'b011100000;
        12'd1265: chroma9 = 9'b011100010;
        12'd1266: chroma9 = 9'b011100100;
        12'd1267: chroma9 = 9'b011100110;
        12'd1268: chroma9 = 9'b011101000;
        12'd1269: chroma9 = 9'b011101010;
        12'd1270: chroma9 = 9'b011101100;
        12'd1271: chroma9 = 9'b011101110;
        12'd1272: chroma9 = 9'b011110000;
        12'd1273: chroma9 = 9'b011110010;
        12'd1274: chroma9 = 9'b011110100;
        12'd1275: chroma9 = 9'b011110110;
        12'd1276: chroma9 = 9'b011111000;
        12'd1277: chroma9 = 9'b011111010;
        12'd1278: chroma9 = 9'b011111100;
        12'd1279: chroma9 = 9'b011111110;
        12'd1280: chroma9 = 9'b100000000;
        12'd1281: chroma9 = 9'b100000010;
        12'd1282: chroma9 = 9'b100000100;
        12'd1283: chroma9 = 9'b100000111;
        12'd1284: chroma9 = 9'b100001001;
        12'd1285: chroma9 = 9'b100001100;
        12'd1286: chroma9 = 9'b100001110;
        12'd1287: chroma9 = 9'b100010001;
        12'd1288: chroma9 = 9'b100010011;
        12'd1289: chroma9 = 9'b100010101;
        12'd1290: chroma9 = 9'b100011000;
        12'd1291: chroma9 = 9'b100011010;
        12'd1292: chroma9 = 9'b100011101;
        12'd1293: chroma9 = 9'b100011111;
        12'd1294: chroma9 = 9'b100100001;
        12'd1295: chroma9 = 9'b100100011;
        12'd1296: chroma9 = 9'b100100110;
        12'd1297: chroma9 = 9'b100101000;
        12'd1298: chroma9 = 9'b100101010;
        12'd1299: chroma9 = 9'b100101100;
        12'd1300: chroma9 = 9'b100101111;
        12'd1301: chroma9 = 9'b100110001;
        12'd1302: chroma9 = 9'b100110011;
        12'd1303: chroma9 = 9'b100110101;
        12'd1304: chroma9 = 9'b100110111;
        12'd1305: chroma9 = 9'b100111001;
        12'd1306: chroma9 = 9'b100111011;
        12'd1307: chroma9 = 9'b100111101;
        12'd1308: chroma9 = 9'b100111111;
        12'd1309: chroma9 = 9'b101000001;
        12'd1310: chroma9 = 9'b101000011;
        12'd1311: chroma9 = 9'b101000100;
        12'd1312: chroma9 = 9'b101000110;
        12'd1313: chroma9 = 9'b101001000;
        12'd1314: chroma9 = 9'b101001010;
        12'd1315: chroma9 = 9'b101001011;
        12'd1316: chroma9 = 9'b101001101;
        12'd1317: chroma9 = 9'b101001110;
        12'd1318: chroma9 = 9'b101010000;
        12'd1319: chroma9 = 9'b101010001;
        12'd1320: chroma9 = 9'b101010011;
        12'd1321: chroma9 = 9'b101010100;
        12'd1322: chroma9 = 9'b101010101;
        12'd1323: chroma9 = 9'b101010111;
        12'd1324: chroma9 = 9'b101011000;
        12'd1325: chroma9 = 9'b101011001;
        12'd1326: chroma9 = 9'b101011010;
        12'd1327: chroma9 = 9'b101011011;
        12'd1328: chroma9 = 9'b101011100;
        12'd1329: chroma9 = 9'b101011101;
        12'd1330: chroma9 = 9'b101011110;
        12'd1331: chroma9 = 9'b101011110;
        12'd1332: chroma9 = 9'b101011111;
        12'd1333: chroma9 = 9'b101100000;
        12'd1334: chroma9 = 9'b101100001;
        12'd1335: chroma9 = 9'b101100001;
        12'd1336: chroma9 = 9'b101100010;
        12'd1337: chroma9 = 9'b101100010;
        12'd1338: chroma9 = 9'b101100010;
        12'd1339: chroma9 = 9'b101100011;
        12'd1340: chroma9 = 9'b101100011;
        12'd1341: chroma9 = 9'b101100011;
        12'd1342: chroma9 = 9'b101100011;
        12'd1343: chroma9 = 9'b101100011;
        12'd1344: chroma9 = 9'b101100011;
        12'd1345: chroma9 = 9'b101100011;
        12'd1346: chroma9 = 9'b101100011;
        12'd1347: chroma9 = 9'b101100011;
        12'd1348: chroma9 = 9'b101100011;
        12'd1349: chroma9 = 9'b101100011;
        12'd1350: chroma9 = 9'b101100010;
        12'd1351: chroma9 = 9'b101100010;
        12'd1352: chroma9 = 9'b101100010;
        12'd1353: chroma9 = 9'b101100001;
        12'd1354: chroma9 = 9'b101100001;
        12'd1355: chroma9 = 9'b101100000;
        12'd1356: chroma9 = 9'b101011111;
        12'd1357: chroma9 = 9'b101011110;
        12'd1358: chroma9 = 9'b101011110;
        12'd1359: chroma9 = 9'b101011101;
        12'd1360: chroma9 = 9'b101011100;
        12'd1361: chroma9 = 9'b101011011;
        12'd1362: chroma9 = 9'b101011010;
        12'd1363: chroma9 = 9'b101011001;
        12'd1364: chroma9 = 9'b101011000;
        12'd1365: chroma9 = 9'b101010111;
        12'd1366: chroma9 = 9'b101010101;
        12'd1367: chroma9 = 9'b101010100;
        12'd1368: chroma9 = 9'b101010011;
        12'd1369: chroma9 = 9'b101010001;
        12'd1370: chroma9 = 9'b101010000;
        12'd1371: chroma9 = 9'b101001110;
        12'd1372: chroma9 = 9'b101001101;
        12'd1373: chroma9 = 9'b101001011;
        12'd1374: chroma9 = 9'b101001010;
        12'd1375: chroma9 = 9'b101001000;
        12'd1376: chroma9 = 9'b101000110;
        12'd1377: chroma9 = 9'b101000100;
        12'd1378: chroma9 = 9'b101000011;
        12'd1379: chroma9 = 9'b101000001;
        12'd1380: chroma9 = 9'b100111111;
        12'd1381: chroma9 = 9'b100111101;
        12'd1382: chroma9 = 9'b100111011;
        12'd1383: chroma9 = 9'b100111001;
        12'd1384: chroma9 = 9'b100110111;
        12'd1385: chroma9 = 9'b100110101;
        12'd1386: chroma9 = 9'b100110011;
        12'd1387: chroma9 = 9'b100110001;
        12'd1388: chroma9 = 9'b100101111;
        12'd1389: chroma9 = 9'b100101100;
        12'd1390: chroma9 = 9'b100101010;
        12'd1391: chroma9 = 9'b100101000;
        12'd1392: chroma9 = 9'b100100110;
        12'd1393: chroma9 = 9'b100100011;
        12'd1394: chroma9 = 9'b100100001;
        12'd1395: chroma9 = 9'b100011111;
        12'd1396: chroma9 = 9'b100011101;
        12'd1397: chroma9 = 9'b100011010;
        12'd1398: chroma9 = 9'b100011000;
        12'd1399: chroma9 = 9'b100010101;
        12'd1400: chroma9 = 9'b100010011;
        12'd1401: chroma9 = 9'b100010001;
        12'd1402: chroma9 = 9'b100001110;
        12'd1403: chroma9 = 9'b100001100;
        12'd1404: chroma9 = 9'b100001001;
        12'd1405: chroma9 = 9'b100000111;
        12'd1406: chroma9 = 9'b100000100;
        12'd1407: chroma9 = 9'b100000010;
        12'd1408: chroma9 = 9'b100000000;
        12'd1409: chroma9 = 9'b011111110;
        12'd1410: chroma9 = 9'b011111100;
        12'd1411: chroma9 = 9'b011111001;
        12'd1412: chroma9 = 9'b011110111;
        12'd1413: chroma9 = 9'b011110100;
        12'd1414: chroma9 = 9'b011110010;
        12'd1415: chroma9 = 9'b011101111;
        12'd1416: chroma9 = 9'b011101101;
        12'd1417: chroma9 = 9'b011101011;
        12'd1418: chroma9 = 9'b011101000;
        12'd1419: chroma9 = 9'b011100110;
        12'd1420: chroma9 = 9'b011100011;
        12'd1421: chroma9 = 9'b011100001;
        12'd1422: chroma9 = 9'b011011111;
        12'd1423: chroma9 = 9'b011011101;
        12'd1424: chroma9 = 9'b011011010;
        12'd1425: chroma9 = 9'b011011000;
        12'd1426: chroma9 = 9'b011010110;
        12'd1427: chroma9 = 9'b011010100;
        12'd1428: chroma9 = 9'b011010001;
        12'd1429: chroma9 = 9'b011001111;
        12'd1430: chroma9 = 9'b011001101;
        12'd1431: chroma9 = 9'b011001011;
        12'd1432: chroma9 = 9'b011001001;
        12'd1433: chroma9 = 9'b011000111;
        12'd1434: chroma9 = 9'b011000101;
        12'd1435: chroma9 = 9'b011000011;
        12'd1436: chroma9 = 9'b011000001;
        12'd1437: chroma9 = 9'b010111111;
        12'd1438: chroma9 = 9'b010111101;
        12'd1439: chroma9 = 9'b010111100;
        12'd1440: chroma9 = 9'b010111010;
        12'd1441: chroma9 = 9'b010111000;
        12'd1442: chroma9 = 9'b010110110;
        12'd1443: chroma9 = 9'b010110101;
        12'd1444: chroma9 = 9'b010110011;
        12'd1445: chroma9 = 9'b010110010;
        12'd1446: chroma9 = 9'b010110000;
        12'd1447: chroma9 = 9'b010101111;
        12'd1448: chroma9 = 9'b010101101;
        12'd1449: chroma9 = 9'b010101100;
        12'd1450: chroma9 = 9'b010101011;
        12'd1451: chroma9 = 9'b010101001;
        12'd1452: chroma9 = 9'b010101000;
        12'd1453: chroma9 = 9'b010100111;
        12'd1454: chroma9 = 9'b010100110;
        12'd1455: chroma9 = 9'b010100101;
        12'd1456: chroma9 = 9'b010100100;
        12'd1457: chroma9 = 9'b010100011;
        12'd1458: chroma9 = 9'b010100010;
        12'd1459: chroma9 = 9'b010100010;
        12'd1460: chroma9 = 9'b010100001;
        12'd1461: chroma9 = 9'b010100000;
        12'd1462: chroma9 = 9'b010011111;
        12'd1463: chroma9 = 9'b010011111;
        12'd1464: chroma9 = 9'b010011110;
        12'd1465: chroma9 = 9'b010011110;
        12'd1466: chroma9 = 9'b010011110;
        12'd1467: chroma9 = 9'b010011101;
        12'd1468: chroma9 = 9'b010011101;
        12'd1469: chroma9 = 9'b010011101;
        12'd1470: chroma9 = 9'b010011101;
        12'd1471: chroma9 = 9'b010011101;
        12'd1472: chroma9 = 9'b010011101;
        12'd1473: chroma9 = 9'b010011101;
        12'd1474: chroma9 = 9'b010011101;
        12'd1475: chroma9 = 9'b010011101;
        12'd1476: chroma9 = 9'b010011101;
        12'd1477: chroma9 = 9'b010011101;
        12'd1478: chroma9 = 9'b010011110;
        12'd1479: chroma9 = 9'b010011110;
        12'd1480: chroma9 = 9'b010011110;
        12'd1481: chroma9 = 9'b010011111;
        12'd1482: chroma9 = 9'b010011111;
        12'd1483: chroma9 = 9'b010100000;
        12'd1484: chroma9 = 9'b010100001;
        12'd1485: chroma9 = 9'b010100010;
        12'd1486: chroma9 = 9'b010100010;
        12'd1487: chroma9 = 9'b010100011;
        12'd1488: chroma9 = 9'b010100100;
        12'd1489: chroma9 = 9'b010100101;
        12'd1490: chroma9 = 9'b010100110;
        12'd1491: chroma9 = 9'b010100111;
        12'd1492: chroma9 = 9'b010101000;
        12'd1493: chroma9 = 9'b010101001;
        12'd1494: chroma9 = 9'b010101011;
        12'd1495: chroma9 = 9'b010101100;
        12'd1496: chroma9 = 9'b010101101;
        12'd1497: chroma9 = 9'b010101111;
        12'd1498: chroma9 = 9'b010110000;
        12'd1499: chroma9 = 9'b010110010;
        12'd1500: chroma9 = 9'b010110011;
        12'd1501: chroma9 = 9'b010110101;
        12'd1502: chroma9 = 9'b010110110;
        12'd1503: chroma9 = 9'b010111000;
        12'd1504: chroma9 = 9'b010111010;
        12'd1505: chroma9 = 9'b010111100;
        12'd1506: chroma9 = 9'b010111101;
        12'd1507: chroma9 = 9'b010111111;
        12'd1508: chroma9 = 9'b011000001;
        12'd1509: chroma9 = 9'b011000011;
        12'd1510: chroma9 = 9'b011000101;
        12'd1511: chroma9 = 9'b011000111;
        12'd1512: chroma9 = 9'b011001001;
        12'd1513: chroma9 = 9'b011001011;
        12'd1514: chroma9 = 9'b011001101;
        12'd1515: chroma9 = 9'b011001111;
        12'd1516: chroma9 = 9'b011010001;
        12'd1517: chroma9 = 9'b011010100;
        12'd1518: chroma9 = 9'b011010110;
        12'd1519: chroma9 = 9'b011011000;
        12'd1520: chroma9 = 9'b011011010;
        12'd1521: chroma9 = 9'b011011101;
        12'd1522: chroma9 = 9'b011011111;
        12'd1523: chroma9 = 9'b011100001;
        12'd1524: chroma9 = 9'b011100011;
        12'd1525: chroma9 = 9'b011100110;
        12'd1526: chroma9 = 9'b011101000;
        12'd1527: chroma9 = 9'b011101011;
        12'd1528: chroma9 = 9'b011101101;
        12'd1529: chroma9 = 9'b011101111;
        12'd1530: chroma9 = 9'b011110010;
        12'd1531: chroma9 = 9'b011110100;
        12'd1532: chroma9 = 9'b011110111;
        12'd1533: chroma9 = 9'b011111001;
        12'd1534: chroma9 = 9'b011111100;
        12'd1535: chroma9 = 9'b011111110;
        12'd1536: chroma9 = 9'b100000000;
        12'd1537: chroma9 = 9'b100000010;
        12'd1538: chroma9 = 9'b100000101;
        12'd1539: chroma9 = 9'b100001000;
        12'd1540: chroma9 = 9'b100001011;
        12'd1541: chroma9 = 9'b100001110;
        12'd1542: chroma9 = 9'b100010000;
        12'd1543: chroma9 = 9'b100010011;
        12'd1544: chroma9 = 9'b100010110;
        12'd1545: chroma9 = 9'b100011001;
        12'd1546: chroma9 = 9'b100011011;
        12'd1547: chroma9 = 9'b100011110;
        12'd1548: chroma9 = 9'b100100001;
        12'd1549: chroma9 = 9'b100100100;
        12'd1550: chroma9 = 9'b100100110;
        12'd1551: chroma9 = 9'b100101001;
        12'd1552: chroma9 = 9'b100101100;
        12'd1553: chroma9 = 9'b100101110;
        12'd1554: chroma9 = 9'b100110001;
        12'd1555: chroma9 = 9'b100110011;
        12'd1556: chroma9 = 9'b100110110;
        12'd1557: chroma9 = 9'b100111000;
        12'd1558: chroma9 = 9'b100111011;
        12'd1559: chroma9 = 9'b100111101;
        12'd1560: chroma9 = 9'b100111111;
        12'd1561: chroma9 = 9'b101000010;
        12'd1562: chroma9 = 9'b101000100;
        12'd1563: chroma9 = 9'b101000110;
        12'd1564: chroma9 = 9'b101001000;
        12'd1565: chroma9 = 9'b101001011;
        12'd1566: chroma9 = 9'b101001101;
        12'd1567: chroma9 = 9'b101001111;
        12'd1568: chroma9 = 9'b101010001;
        12'd1569: chroma9 = 9'b101010011;
        12'd1570: chroma9 = 9'b101010101;
        12'd1571: chroma9 = 9'b101010111;
        12'd1572: chroma9 = 9'b101011000;
        12'd1573: chroma9 = 9'b101011010;
        12'd1574: chroma9 = 9'b101011100;
        12'd1575: chroma9 = 9'b101011110;
        12'd1576: chroma9 = 9'b101011111;
        12'd1577: chroma9 = 9'b101100001;
        12'd1578: chroma9 = 9'b101100010;
        12'd1579: chroma9 = 9'b101100100;
        12'd1580: chroma9 = 9'b101100101;
        12'd1581: chroma9 = 9'b101100110;
        12'd1582: chroma9 = 9'b101100111;
        12'd1583: chroma9 = 9'b101101001;
        12'd1584: chroma9 = 9'b101101010;
        12'd1585: chroma9 = 9'b101101011;
        12'd1586: chroma9 = 9'b101101100;
        12'd1587: chroma9 = 9'b101101101;
        12'd1588: chroma9 = 9'b101101110;
        12'd1589: chroma9 = 9'b101101110;
        12'd1590: chroma9 = 9'b101101111;
        12'd1591: chroma9 = 9'b101110000;
        12'd1592: chroma9 = 9'b101110000;
        12'd1593: chroma9 = 9'b101110001;
        12'd1594: chroma9 = 9'b101110001;
        12'd1595: chroma9 = 9'b101110010;
        12'd1596: chroma9 = 9'b101110010;
        12'd1597: chroma9 = 9'b101110010;
        12'd1598: chroma9 = 9'b101110010;
        12'd1599: chroma9 = 9'b101110010;
        12'd1600: chroma9 = 9'b101110010;
        12'd1601: chroma9 = 9'b101110010;
        12'd1602: chroma9 = 9'b101110010;
        12'd1603: chroma9 = 9'b101110010;
        12'd1604: chroma9 = 9'b101110010;
        12'd1605: chroma9 = 9'b101110010;
        12'd1606: chroma9 = 9'b101110001;
        12'd1607: chroma9 = 9'b101110001;
        12'd1608: chroma9 = 9'b101110000;
        12'd1609: chroma9 = 9'b101110000;
        12'd1610: chroma9 = 9'b101101111;
        12'd1611: chroma9 = 9'b101101110;
        12'd1612: chroma9 = 9'b101101110;
        12'd1613: chroma9 = 9'b101101101;
        12'd1614: chroma9 = 9'b101101100;
        12'd1615: chroma9 = 9'b101101011;
        12'd1616: chroma9 = 9'b101101010;
        12'd1617: chroma9 = 9'b101101001;
        12'd1618: chroma9 = 9'b101100111;
        12'd1619: chroma9 = 9'b101100110;
        12'd1620: chroma9 = 9'b101100101;
        12'd1621: chroma9 = 9'b101100100;
        12'd1622: chroma9 = 9'b101100010;
        12'd1623: chroma9 = 9'b101100001;
        12'd1624: chroma9 = 9'b101011111;
        12'd1625: chroma9 = 9'b101011110;
        12'd1626: chroma9 = 9'b101011100;
        12'd1627: chroma9 = 9'b101011010;
        12'd1628: chroma9 = 9'b101011000;
        12'd1629: chroma9 = 9'b101010111;
        12'd1630: chroma9 = 9'b101010101;
        12'd1631: chroma9 = 9'b101010011;
        12'd1632: chroma9 = 9'b101010001;
        12'd1633: chroma9 = 9'b101001111;
        12'd1634: chroma9 = 9'b101001101;
        12'd1635: chroma9 = 9'b101001011;
        12'd1636: chroma9 = 9'b101001000;
        12'd1637: chroma9 = 9'b101000110;
        12'd1638: chroma9 = 9'b101000100;
        12'd1639: chroma9 = 9'b101000010;
        12'd1640: chroma9 = 9'b100111111;
        12'd1641: chroma9 = 9'b100111101;
        12'd1642: chroma9 = 9'b100111011;
        12'd1643: chroma9 = 9'b100111000;
        12'd1644: chroma9 = 9'b100110110;
        12'd1645: chroma9 = 9'b100110011;
        12'd1646: chroma9 = 9'b100110001;
        12'd1647: chroma9 = 9'b100101110;
        12'd1648: chroma9 = 9'b100101100;
        12'd1649: chroma9 = 9'b100101001;
        12'd1650: chroma9 = 9'b100100110;
        12'd1651: chroma9 = 9'b100100100;
        12'd1652: chroma9 = 9'b100100001;
        12'd1653: chroma9 = 9'b100011110;
        12'd1654: chroma9 = 9'b100011011;
        12'd1655: chroma9 = 9'b100011001;
        12'd1656: chroma9 = 9'b100010110;
        12'd1657: chroma9 = 9'b100010011;
        12'd1658: chroma9 = 9'b100010000;
        12'd1659: chroma9 = 9'b100001110;
        12'd1660: chroma9 = 9'b100001011;
        12'd1661: chroma9 = 9'b100001000;
        12'd1662: chroma9 = 9'b100000101;
        12'd1663: chroma9 = 9'b100000010;
        12'd1664: chroma9 = 9'b100000000;
        12'd1665: chroma9 = 9'b011111110;
        12'd1666: chroma9 = 9'b011111011;
        12'd1667: chroma9 = 9'b011111000;
        12'd1668: chroma9 = 9'b011110101;
        12'd1669: chroma9 = 9'b011110010;
        12'd1670: chroma9 = 9'b011110000;
        12'd1671: chroma9 = 9'b011101101;
        12'd1672: chroma9 = 9'b011101010;
        12'd1673: chroma9 = 9'b011100111;
        12'd1674: chroma9 = 9'b011100101;
        12'd1675: chroma9 = 9'b011100010;
        12'd1676: chroma9 = 9'b011011111;
        12'd1677: chroma9 = 9'b011011100;
        12'd1678: chroma9 = 9'b011011010;
        12'd1679: chroma9 = 9'b011010111;
        12'd1680: chroma9 = 9'b011010100;
        12'd1681: chroma9 = 9'b011010010;
        12'd1682: chroma9 = 9'b011001111;
        12'd1683: chroma9 = 9'b011001101;
        12'd1684: chroma9 = 9'b011001010;
        12'd1685: chroma9 = 9'b011001000;
        12'd1686: chroma9 = 9'b011000101;
        12'd1687: chroma9 = 9'b011000011;
        12'd1688: chroma9 = 9'b011000001;
        12'd1689: chroma9 = 9'b010111110;
        12'd1690: chroma9 = 9'b010111100;
        12'd1691: chroma9 = 9'b010111010;
        12'd1692: chroma9 = 9'b010111000;
        12'd1693: chroma9 = 9'b010110101;
        12'd1694: chroma9 = 9'b010110011;
        12'd1695: chroma9 = 9'b010110001;
        12'd1696: chroma9 = 9'b010101111;
        12'd1697: chroma9 = 9'b010101101;
        12'd1698: chroma9 = 9'b010101011;
        12'd1699: chroma9 = 9'b010101001;
        12'd1700: chroma9 = 9'b010101000;
        12'd1701: chroma9 = 9'b010100110;
        12'd1702: chroma9 = 9'b010100100;
        12'd1703: chroma9 = 9'b010100010;
        12'd1704: chroma9 = 9'b010100001;
        12'd1705: chroma9 = 9'b010011111;
        12'd1706: chroma9 = 9'b010011110;
        12'd1707: chroma9 = 9'b010011100;
        12'd1708: chroma9 = 9'b010011011;
        12'd1709: chroma9 = 9'b010011010;
        12'd1710: chroma9 = 9'b010011001;
        12'd1711: chroma9 = 9'b010010111;
        12'd1712: chroma9 = 9'b010010110;
        12'd1713: chroma9 = 9'b010010101;
        12'd1714: chroma9 = 9'b010010100;
        12'd1715: chroma9 = 9'b010010011;
        12'd1716: chroma9 = 9'b010010010;
        12'd1717: chroma9 = 9'b010010010;
        12'd1718: chroma9 = 9'b010010001;
        12'd1719: chroma9 = 9'b010010000;
        12'd1720: chroma9 = 9'b010010000;
        12'd1721: chroma9 = 9'b010001111;
        12'd1722: chroma9 = 9'b010001111;
        12'd1723: chroma9 = 9'b010001110;
        12'd1724: chroma9 = 9'b010001110;
        12'd1725: chroma9 = 9'b010001110;
        12'd1726: chroma9 = 9'b010001110;
        12'd1727: chroma9 = 9'b010001110;
        12'd1728: chroma9 = 9'b010001110;
        12'd1729: chroma9 = 9'b010001110;
        12'd1730: chroma9 = 9'b010001110;
        12'd1731: chroma9 = 9'b010001110;
        12'd1732: chroma9 = 9'b010001110;
        12'd1733: chroma9 = 9'b010001110;
        12'd1734: chroma9 = 9'b010001111;
        12'd1735: chroma9 = 9'b010001111;
        12'd1736: chroma9 = 9'b010010000;
        12'd1737: chroma9 = 9'b010010000;
        12'd1738: chroma9 = 9'b010010001;
        12'd1739: chroma9 = 9'b010010010;
        12'd1740: chroma9 = 9'b010010010;
        12'd1741: chroma9 = 9'b010010011;
        12'd1742: chroma9 = 9'b010010100;
        12'd1743: chroma9 = 9'b010010101;
        12'd1744: chroma9 = 9'b010010110;
        12'd1745: chroma9 = 9'b010010111;
        12'd1746: chroma9 = 9'b010011001;
        12'd1747: chroma9 = 9'b010011010;
        12'd1748: chroma9 = 9'b010011011;
        12'd1749: chroma9 = 9'b010011100;
        12'd1750: chroma9 = 9'b010011110;
        12'd1751: chroma9 = 9'b010011111;
        12'd1752: chroma9 = 9'b010100001;
        12'd1753: chroma9 = 9'b010100010;
        12'd1754: chroma9 = 9'b010100100;
        12'd1755: chroma9 = 9'b010100110;
        12'd1756: chroma9 = 9'b010101000;
        12'd1757: chroma9 = 9'b010101001;
        12'd1758: chroma9 = 9'b010101011;
        12'd1759: chroma9 = 9'b010101101;
        12'd1760: chroma9 = 9'b010101111;
        12'd1761: chroma9 = 9'b010110001;
        12'd1762: chroma9 = 9'b010110011;
        12'd1763: chroma9 = 9'b010110101;
        12'd1764: chroma9 = 9'b010111000;
        12'd1765: chroma9 = 9'b010111010;
        12'd1766: chroma9 = 9'b010111100;
        12'd1767: chroma9 = 9'b010111110;
        12'd1768: chroma9 = 9'b011000001;
        12'd1769: chroma9 = 9'b011000011;
        12'd1770: chroma9 = 9'b011000101;
        12'd1771: chroma9 = 9'b011001000;
        12'd1772: chroma9 = 9'b011001010;
        12'd1773: chroma9 = 9'b011001101;
        12'd1774: chroma9 = 9'b011001111;
        12'd1775: chroma9 = 9'b011010010;
        12'd1776: chroma9 = 9'b011010100;
        12'd1777: chroma9 = 9'b011010111;
        12'd1778: chroma9 = 9'b011011010;
        12'd1779: chroma9 = 9'b011011100;
        12'd1780: chroma9 = 9'b011011111;
        12'd1781: chroma9 = 9'b011100010;
        12'd1782: chroma9 = 9'b011100101;
        12'd1783: chroma9 = 9'b011100111;
        12'd1784: chroma9 = 9'b011101010;
        12'd1785: chroma9 = 9'b011101101;
        12'd1786: chroma9 = 9'b011110000;
        12'd1787: chroma9 = 9'b011110010;
        12'd1788: chroma9 = 9'b011110101;
        12'd1789: chroma9 = 9'b011111000;
        12'd1790: chroma9 = 9'b011111011;
        12'd1791: chroma9 = 9'b011111110;
        12'd1792: chroma9 = 9'b100000000;
        12'd1793: chroma9 = 9'b100000011;
        12'd1794: chroma9 = 9'b100000110;
        12'd1795: chroma9 = 9'b100001001;
        12'd1796: chroma9 = 9'b100001100;
        12'd1797: chroma9 = 9'b100001111;
        12'd1798: chroma9 = 9'b100010011;
        12'd1799: chroma9 = 9'b100010110;
        12'd1800: chroma9 = 9'b100011001;
        12'd1801: chroma9 = 9'b100011100;
        12'd1802: chroma9 = 9'b100011111;
        12'd1803: chroma9 = 9'b100100010;
        12'd1804: chroma9 = 9'b100100101;
        12'd1805: chroma9 = 9'b100101000;
        12'd1806: chroma9 = 9'b100101011;
        12'd1807: chroma9 = 9'b100101110;
        12'd1808: chroma9 = 9'b100110001;
        12'd1809: chroma9 = 9'b100110100;
        12'd1810: chroma9 = 9'b100110111;
        12'd1811: chroma9 = 9'b100111010;
        12'd1812: chroma9 = 9'b100111101;
        12'd1813: chroma9 = 9'b101000000;
        12'd1814: chroma9 = 9'b101000010;
        12'd1815: chroma9 = 9'b101000101;
        12'd1816: chroma9 = 9'b101001000;
        12'd1817: chroma9 = 9'b101001010;
        12'd1818: chroma9 = 9'b101001101;
        12'd1819: chroma9 = 9'b101001111;
        12'd1820: chroma9 = 9'b101010010;
        12'd1821: chroma9 = 9'b101010100;
        12'd1822: chroma9 = 9'b101010111;
        12'd1823: chroma9 = 9'b101011001;
        12'd1824: chroma9 = 9'b101011011;
        12'd1825: chroma9 = 9'b101011110;
        12'd1826: chroma9 = 9'b101100000;
        12'd1827: chroma9 = 9'b101100010;
        12'd1828: chroma9 = 9'b101100100;
        12'd1829: chroma9 = 9'b101100110;
        12'd1830: chroma9 = 9'b101101000;
        12'd1831: chroma9 = 9'b101101010;
        12'd1832: chroma9 = 9'b101101100;
        12'd1833: chroma9 = 9'b101101101;
        12'd1834: chroma9 = 9'b101101111;
        12'd1835: chroma9 = 9'b101110001;
        12'd1836: chroma9 = 9'b101110010;
        12'd1837: chroma9 = 9'b101110100;
        12'd1838: chroma9 = 9'b101110101;
        12'd1839: chroma9 = 9'b101110110;
        12'd1840: chroma9 = 9'b101111000;
        12'd1841: chroma9 = 9'b101111001;
        12'd1842: chroma9 = 9'b101111010;
        12'd1843: chroma9 = 9'b101111011;
        12'd1844: chroma9 = 9'b101111100;
        12'd1845: chroma9 = 9'b101111101;
        12'd1846: chroma9 = 9'b101111110;
        12'd1847: chroma9 = 9'b101111110;
        12'd1848: chroma9 = 9'b101111111;
        12'd1849: chroma9 = 9'b110000000;
        12'd1850: chroma9 = 9'b110000000;
        12'd1851: chroma9 = 9'b110000001;
        12'd1852: chroma9 = 9'b110000001;
        12'd1853: chroma9 = 9'b110000001;
        12'd1854: chroma9 = 9'b110000001;
        12'd1855: chroma9 = 9'b110000001;
        12'd1856: chroma9 = 9'b110000001;
        12'd1857: chroma9 = 9'b110000001;
        12'd1858: chroma9 = 9'b110000001;
        12'd1859: chroma9 = 9'b110000001;
        12'd1860: chroma9 = 9'b110000001;
        12'd1861: chroma9 = 9'b110000001;
        12'd1862: chroma9 = 9'b110000000;
        12'd1863: chroma9 = 9'b110000000;
        12'd1864: chroma9 = 9'b101111111;
        12'd1865: chroma9 = 9'b101111110;
        12'd1866: chroma9 = 9'b101111110;
        12'd1867: chroma9 = 9'b101111101;
        12'd1868: chroma9 = 9'b101111100;
        12'd1869: chroma9 = 9'b101111011;
        12'd1870: chroma9 = 9'b101111010;
        12'd1871: chroma9 = 9'b101111001;
        12'd1872: chroma9 = 9'b101111000;
        12'd1873: chroma9 = 9'b101110110;
        12'd1874: chroma9 = 9'b101110101;
        12'd1875: chroma9 = 9'b101110100;
        12'd1876: chroma9 = 9'b101110010;
        12'd1877: chroma9 = 9'b101110001;
        12'd1878: chroma9 = 9'b101101111;
        12'd1879: chroma9 = 9'b101101101;
        12'd1880: chroma9 = 9'b101101100;
        12'd1881: chroma9 = 9'b101101010;
        12'd1882: chroma9 = 9'b101101000;
        12'd1883: chroma9 = 9'b101100110;
        12'd1884: chroma9 = 9'b101100100;
        12'd1885: chroma9 = 9'b101100010;
        12'd1886: chroma9 = 9'b101100000;
        12'd1887: chroma9 = 9'b101011110;
        12'd1888: chroma9 = 9'b101011011;
        12'd1889: chroma9 = 9'b101011001;
        12'd1890: chroma9 = 9'b101010111;
        12'd1891: chroma9 = 9'b101010100;
        12'd1892: chroma9 = 9'b101010010;
        12'd1893: chroma9 = 9'b101001111;
        12'd1894: chroma9 = 9'b101001101;
        12'd1895: chroma9 = 9'b101001010;
        12'd1896: chroma9 = 9'b101001000;
        12'd1897: chroma9 = 9'b101000101;
        12'd1898: chroma9 = 9'b101000010;
        12'd1899: chroma9 = 9'b101000000;
        12'd1900: chroma9 = 9'b100111101;
        12'd1901: chroma9 = 9'b100111010;
        12'd1902: chroma9 = 9'b100110111;
        12'd1903: chroma9 = 9'b100110100;
        12'd1904: chroma9 = 9'b100110001;
        12'd1905: chroma9 = 9'b100101110;
        12'd1906: chroma9 = 9'b100101011;
        12'd1907: chroma9 = 9'b100101000;
        12'd1908: chroma9 = 9'b100100101;
        12'd1909: chroma9 = 9'b100100010;
        12'd1910: chroma9 = 9'b100011111;
        12'd1911: chroma9 = 9'b100011100;
        12'd1912: chroma9 = 9'b100011001;
        12'd1913: chroma9 = 9'b100010110;
        12'd1914: chroma9 = 9'b100010011;
        12'd1915: chroma9 = 9'b100001111;
        12'd1916: chroma9 = 9'b100001100;
        12'd1917: chroma9 = 9'b100001001;
        12'd1918: chroma9 = 9'b100000110;
        12'd1919: chroma9 = 9'b100000011;
        12'd1920: chroma9 = 9'b100000000;
        12'd1921: chroma9 = 9'b011111101;
        12'd1922: chroma9 = 9'b011111010;
        12'd1923: chroma9 = 9'b011110111;
        12'd1924: chroma9 = 9'b011110100;
        12'd1925: chroma9 = 9'b011110001;
        12'd1926: chroma9 = 9'b011101101;
        12'd1927: chroma9 = 9'b011101010;
        12'd1928: chroma9 = 9'b011100111;
        12'd1929: chroma9 = 9'b011100100;
        12'd1930: chroma9 = 9'b011100001;
        12'd1931: chroma9 = 9'b011011110;
        12'd1932: chroma9 = 9'b011011011;
        12'd1933: chroma9 = 9'b011011000;
        12'd1934: chroma9 = 9'b011010101;
        12'd1935: chroma9 = 9'b011010010;
        12'd1936: chroma9 = 9'b011001111;
        12'd1937: chroma9 = 9'b011001100;
        12'd1938: chroma9 = 9'b011001001;
        12'd1939: chroma9 = 9'b011000110;
        12'd1940: chroma9 = 9'b011000011;
        12'd1941: chroma9 = 9'b011000000;
        12'd1942: chroma9 = 9'b010111110;
        12'd1943: chroma9 = 9'b010111011;
        12'd1944: chroma9 = 9'b010111000;
        12'd1945: chroma9 = 9'b010110110;
        12'd1946: chroma9 = 9'b010110011;
        12'd1947: chroma9 = 9'b010110001;
        12'd1948: chroma9 = 9'b010101110;
        12'd1949: chroma9 = 9'b010101100;
        12'd1950: chroma9 = 9'b010101001;
        12'd1951: chroma9 = 9'b010100111;
        12'd1952: chroma9 = 9'b010100101;
        12'd1953: chroma9 = 9'b010100010;
        12'd1954: chroma9 = 9'b010100000;
        12'd1955: chroma9 = 9'b010011110;
        12'd1956: chroma9 = 9'b010011100;
        12'd1957: chroma9 = 9'b010011010;
        12'd1958: chroma9 = 9'b010011000;
        12'd1959: chroma9 = 9'b010010110;
        12'd1960: chroma9 = 9'b010010100;
        12'd1961: chroma9 = 9'b010010011;
        12'd1962: chroma9 = 9'b010010001;
        12'd1963: chroma9 = 9'b010001111;
        12'd1964: chroma9 = 9'b010001110;
        12'd1965: chroma9 = 9'b010001100;
        12'd1966: chroma9 = 9'b010001011;
        12'd1967: chroma9 = 9'b010001010;
        12'd1968: chroma9 = 9'b010001000;
        12'd1969: chroma9 = 9'b010000111;
        12'd1970: chroma9 = 9'b010000110;
        12'd1971: chroma9 = 9'b010000101;
        12'd1972: chroma9 = 9'b010000100;
        12'd1973: chroma9 = 9'b010000011;
        12'd1974: chroma9 = 9'b010000010;
        12'd1975: chroma9 = 9'b010000010;
        12'd1976: chroma9 = 9'b010000001;
        12'd1977: chroma9 = 9'b010000000;
        12'd1978: chroma9 = 9'b010000000;
        12'd1979: chroma9 = 9'b001111111;
        12'd1980: chroma9 = 9'b001111111;
        12'd1981: chroma9 = 9'b001111111;
        12'd1982: chroma9 = 9'b001111111;
        12'd1983: chroma9 = 9'b001111111;
        12'd1984: chroma9 = 9'b001111111;
        12'd1985: chroma9 = 9'b001111111;
        12'd1986: chroma9 = 9'b001111111;
        12'd1987: chroma9 = 9'b001111111;
        12'd1988: chroma9 = 9'b001111111;
        12'd1989: chroma9 = 9'b001111111;
        12'd1990: chroma9 = 9'b010000000;
        12'd1991: chroma9 = 9'b010000000;
        12'd1992: chroma9 = 9'b010000001;
        12'd1993: chroma9 = 9'b010000010;
        12'd1994: chroma9 = 9'b010000010;
        12'd1995: chroma9 = 9'b010000011;
        12'd1996: chroma9 = 9'b010000100;
        12'd1997: chroma9 = 9'b010000101;
        12'd1998: chroma9 = 9'b010000110;
        12'd1999: chroma9 = 9'b010000111;
        12'd2000: chroma9 = 9'b010001000;
        12'd2001: chroma9 = 9'b010001010;
        12'd2002: chroma9 = 9'b010001011;
        12'd2003: chroma9 = 9'b010001100;
        12'd2004: chroma9 = 9'b010001110;
        12'd2005: chroma9 = 9'b010001111;
        12'd2006: chroma9 = 9'b010010001;
        12'd2007: chroma9 = 9'b010010011;
        12'd2008: chroma9 = 9'b010010100;
        12'd2009: chroma9 = 9'b010010110;
        12'd2010: chroma9 = 9'b010011000;
        12'd2011: chroma9 = 9'b010011010;
        12'd2012: chroma9 = 9'b010011100;
        12'd2013: chroma9 = 9'b010011110;
        12'd2014: chroma9 = 9'b010100000;
        12'd2015: chroma9 = 9'b010100010;
        12'd2016: chroma9 = 9'b010100101;
        12'd2017: chroma9 = 9'b010100111;
        12'd2018: chroma9 = 9'b010101001;
        12'd2019: chroma9 = 9'b010101100;
        12'd2020: chroma9 = 9'b010101110;
        12'd2021: chroma9 = 9'b010110001;
        12'd2022: chroma9 = 9'b010110011;
        12'd2023: chroma9 = 9'b010110110;
        12'd2024: chroma9 = 9'b010111000;
        12'd2025: chroma9 = 9'b010111011;
        12'd2026: chroma9 = 9'b010111110;
        12'd2027: chroma9 = 9'b011000000;
        12'd2028: chroma9 = 9'b011000011;
        12'd2029: chroma9 = 9'b011000110;
        12'd2030: chroma9 = 9'b011001001;
        12'd2031: chroma9 = 9'b011001100;
        12'd2032: chroma9 = 9'b011001111;
        12'd2033: chroma9 = 9'b011010010;
        12'd2034: chroma9 = 9'b011010101;
        12'd2035: chroma9 = 9'b011011000;
        12'd2036: chroma9 = 9'b011011011;
        12'd2037: chroma9 = 9'b011011110;
        12'd2038: chroma9 = 9'b011100001;
        12'd2039: chroma9 = 9'b011100100;
        12'd2040: chroma9 = 9'b011100111;
        12'd2041: chroma9 = 9'b011101010;
        12'd2042: chroma9 = 9'b011101101;
        12'd2043: chroma9 = 9'b011110001;
        12'd2044: chroma9 = 9'b011110100;
        12'd2045: chroma9 = 9'b011110111;
        12'd2046: chroma9 = 9'b011111010;
        12'd2047: chroma9 = 9'b011111101;
        12'd2048: chroma9 = 9'b100000000;
        12'd2049: chroma9 = 9'b100000011;
        12'd2050: chroma9 = 9'b100000111;
        12'd2051: chroma9 = 9'b100001010;
        12'd2052: chroma9 = 9'b100001110;
        12'd2053: chroma9 = 9'b100010001;
        12'd2054: chroma9 = 9'b100010101;
        12'd2055: chroma9 = 9'b100011000;
        12'd2056: chroma9 = 9'b100011100;
        12'd2057: chroma9 = 9'b100011111;
        12'd2058: chroma9 = 9'b100100011;
        12'd2059: chroma9 = 9'b100100110;
        12'd2060: chroma9 = 9'b100101010;
        12'd2061: chroma9 = 9'b100101101;
        12'd2062: chroma9 = 9'b100110000;
        12'd2063: chroma9 = 9'b100110100;
        12'd2064: chroma9 = 9'b100110111;
        12'd2065: chroma9 = 9'b100111010;
        12'd2066: chroma9 = 9'b100111101;
        12'd2067: chroma9 = 9'b101000001;
        12'd2068: chroma9 = 9'b101000100;
        12'd2069: chroma9 = 9'b101000111;
        12'd2070: chroma9 = 9'b101001010;
        12'd2071: chroma9 = 9'b101001101;
        12'd2072: chroma9 = 9'b101010000;
        12'd2073: chroma9 = 9'b101010011;
        12'd2074: chroma9 = 9'b101010110;
        12'd2075: chroma9 = 9'b101011001;
        12'd2076: chroma9 = 9'b101011011;
        12'd2077: chroma9 = 9'b101011110;
        12'd2078: chroma9 = 9'b101100001;
        12'd2079: chroma9 = 9'b101100011;
        12'd2080: chroma9 = 9'b101100110;
        12'd2081: chroma9 = 9'b101101001;
        12'd2082: chroma9 = 9'b101101011;
        12'd2083: chroma9 = 9'b101101101;
        12'd2084: chroma9 = 9'b101110000;
        12'd2085: chroma9 = 9'b101110010;
        12'd2086: chroma9 = 9'b101110100;
        12'd2087: chroma9 = 9'b101110110;
        12'd2088: chroma9 = 9'b101111000;
        12'd2089: chroma9 = 9'b101111010;
        12'd2090: chroma9 = 9'b101111100;
        12'd2091: chroma9 = 9'b101111110;
        12'd2092: chroma9 = 9'b101111111;
        12'd2093: chroma9 = 9'b110000001;
        12'd2094: chroma9 = 9'b110000011;
        12'd2095: chroma9 = 9'b110000100;
        12'd2096: chroma9 = 9'b110000101;
        12'd2097: chroma9 = 9'b110000111;
        12'd2098: chroma9 = 9'b110001000;
        12'd2099: chroma9 = 9'b110001001;
        12'd2100: chroma9 = 9'b110001010;
        12'd2101: chroma9 = 9'b110001011;
        12'd2102: chroma9 = 9'b110001100;
        12'd2103: chroma9 = 9'b110001101;
        12'd2104: chroma9 = 9'b110001110;
        12'd2105: chroma9 = 9'b110001110;
        12'd2106: chroma9 = 9'b110001111;
        12'd2107: chroma9 = 9'b110001111;
        12'd2108: chroma9 = 9'b110010000;
        12'd2109: chroma9 = 9'b110010000;
        12'd2110: chroma9 = 9'b110010000;
        12'd2111: chroma9 = 9'b110010000;
        12'd2112: chroma9 = 9'b110010000;
        12'd2113: chroma9 = 9'b110010000;
        12'd2114: chroma9 = 9'b110010000;
        12'd2115: chroma9 = 9'b110010000;
        12'd2116: chroma9 = 9'b110010000;
        12'd2117: chroma9 = 9'b110001111;
        12'd2118: chroma9 = 9'b110001111;
        12'd2119: chroma9 = 9'b110001110;
        12'd2120: chroma9 = 9'b110001110;
        12'd2121: chroma9 = 9'b110001101;
        12'd2122: chroma9 = 9'b110001100;
        12'd2123: chroma9 = 9'b110001011;
        12'd2124: chroma9 = 9'b110001010;
        12'd2125: chroma9 = 9'b110001001;
        12'd2126: chroma9 = 9'b110001000;
        12'd2127: chroma9 = 9'b110000111;
        12'd2128: chroma9 = 9'b110000101;
        12'd2129: chroma9 = 9'b110000100;
        12'd2130: chroma9 = 9'b110000011;
        12'd2131: chroma9 = 9'b110000001;
        12'd2132: chroma9 = 9'b101111111;
        12'd2133: chroma9 = 9'b101111110;
        12'd2134: chroma9 = 9'b101111100;
        12'd2135: chroma9 = 9'b101111010;
        12'd2136: chroma9 = 9'b101111000;
        12'd2137: chroma9 = 9'b101110110;
        12'd2138: chroma9 = 9'b101110100;
        12'd2139: chroma9 = 9'b101110010;
        12'd2140: chroma9 = 9'b101110000;
        12'd2141: chroma9 = 9'b101101101;
        12'd2142: chroma9 = 9'b101101011;
        12'd2143: chroma9 = 9'b101101001;
        12'd2144: chroma9 = 9'b101100110;
        12'd2145: chroma9 = 9'b101100011;
        12'd2146: chroma9 = 9'b101100001;
        12'd2147: chroma9 = 9'b101011110;
        12'd2148: chroma9 = 9'b101011011;
        12'd2149: chroma9 = 9'b101011001;
        12'd2150: chroma9 = 9'b101010110;
        12'd2151: chroma9 = 9'b101010011;
        12'd2152: chroma9 = 9'b101010000;
        12'd2153: chroma9 = 9'b101001101;
        12'd2154: chroma9 = 9'b101001010;
        12'd2155: chroma9 = 9'b101000111;
        12'd2156: chroma9 = 9'b101000100;
        12'd2157: chroma9 = 9'b101000001;
        12'd2158: chroma9 = 9'b100111101;
        12'd2159: chroma9 = 9'b100111010;
        12'd2160: chroma9 = 9'b100110111;
        12'd2161: chroma9 = 9'b100110100;
        12'd2162: chroma9 = 9'b100110000;
        12'd2163: chroma9 = 9'b100101101;
        12'd2164: chroma9 = 9'b100101010;
        12'd2165: chroma9 = 9'b100100110;
        12'd2166: chroma9 = 9'b100100011;
        12'd2167: chroma9 = 9'b100011111;
        12'd2168: chroma9 = 9'b100011100;
        12'd2169: chroma9 = 9'b100011000;
        12'd2170: chroma9 = 9'b100010101;
        12'd2171: chroma9 = 9'b100010001;
        12'd2172: chroma9 = 9'b100001110;
        12'd2173: chroma9 = 9'b100001010;
        12'd2174: chroma9 = 9'b100000111;
        12'd2175: chroma9 = 9'b100000011;
        12'd2176: chroma9 = 9'b100000000;
        12'd2177: chroma9 = 9'b011111101;
        12'd2178: chroma9 = 9'b011111001;
        12'd2179: chroma9 = 9'b011110110;
        12'd2180: chroma9 = 9'b011110010;
        12'd2181: chroma9 = 9'b011101111;
        12'd2182: chroma9 = 9'b011101011;
        12'd2183: chroma9 = 9'b011101000;
        12'd2184: chroma9 = 9'b011100100;
        12'd2185: chroma9 = 9'b011100001;
        12'd2186: chroma9 = 9'b011011101;
        12'd2187: chroma9 = 9'b011011010;
        12'd2188: chroma9 = 9'b011010110;
        12'd2189: chroma9 = 9'b011010011;
        12'd2190: chroma9 = 9'b011010000;
        12'd2191: chroma9 = 9'b011001100;
        12'd2192: chroma9 = 9'b011001001;
        12'd2193: chroma9 = 9'b011000110;
        12'd2194: chroma9 = 9'b011000011;
        12'd2195: chroma9 = 9'b010111111;
        12'd2196: chroma9 = 9'b010111100;
        12'd2197: chroma9 = 9'b010111001;
        12'd2198: chroma9 = 9'b010110110;
        12'd2199: chroma9 = 9'b010110011;
        12'd2200: chroma9 = 9'b010110000;
        12'd2201: chroma9 = 9'b010101101;
        12'd2202: chroma9 = 9'b010101010;
        12'd2203: chroma9 = 9'b010100111;
        12'd2204: chroma9 = 9'b010100101;
        12'd2205: chroma9 = 9'b010100010;
        12'd2206: chroma9 = 9'b010011111;
        12'd2207: chroma9 = 9'b010011101;
        12'd2208: chroma9 = 9'b010011010;
        12'd2209: chroma9 = 9'b010010111;
        12'd2210: chroma9 = 9'b010010101;
        12'd2211: chroma9 = 9'b010010011;
        12'd2212: chroma9 = 9'b010010000;
        12'd2213: chroma9 = 9'b010001110;
        12'd2214: chroma9 = 9'b010001100;
        12'd2215: chroma9 = 9'b010001010;
        12'd2216: chroma9 = 9'b010001000;
        12'd2217: chroma9 = 9'b010000110;
        12'd2218: chroma9 = 9'b010000100;
        12'd2219: chroma9 = 9'b010000010;
        12'd2220: chroma9 = 9'b010000001;
        12'd2221: chroma9 = 9'b001111111;
        12'd2222: chroma9 = 9'b001111101;
        12'd2223: chroma9 = 9'b001111100;
        12'd2224: chroma9 = 9'b001111011;
        12'd2225: chroma9 = 9'b001111001;
        12'd2226: chroma9 = 9'b001111000;
        12'd2227: chroma9 = 9'b001110111;
        12'd2228: chroma9 = 9'b001110110;
        12'd2229: chroma9 = 9'b001110101;
        12'd2230: chroma9 = 9'b001110100;
        12'd2231: chroma9 = 9'b001110011;
        12'd2232: chroma9 = 9'b001110010;
        12'd2233: chroma9 = 9'b001110010;
        12'd2234: chroma9 = 9'b001110001;
        12'd2235: chroma9 = 9'b001110001;
        12'd2236: chroma9 = 9'b001110000;
        12'd2237: chroma9 = 9'b001110000;
        12'd2238: chroma9 = 9'b001110000;
        12'd2239: chroma9 = 9'b001110000;
        12'd2240: chroma9 = 9'b001110000;
        12'd2241: chroma9 = 9'b001110000;
        12'd2242: chroma9 = 9'b001110000;
        12'd2243: chroma9 = 9'b001110000;
        12'd2244: chroma9 = 9'b001110000;
        12'd2245: chroma9 = 9'b001110001;
        12'd2246: chroma9 = 9'b001110001;
        12'd2247: chroma9 = 9'b001110010;
        12'd2248: chroma9 = 9'b001110010;
        12'd2249: chroma9 = 9'b001110011;
        12'd2250: chroma9 = 9'b001110100;
        12'd2251: chroma9 = 9'b001110101;
        12'd2252: chroma9 = 9'b001110110;
        12'd2253: chroma9 = 9'b001110111;
        12'd2254: chroma9 = 9'b001111000;
        12'd2255: chroma9 = 9'b001111001;
        12'd2256: chroma9 = 9'b001111011;
        12'd2257: chroma9 = 9'b001111100;
        12'd2258: chroma9 = 9'b001111101;
        12'd2259: chroma9 = 9'b001111111;
        12'd2260: chroma9 = 9'b010000001;
        12'd2261: chroma9 = 9'b010000010;
        12'd2262: chroma9 = 9'b010000100;
        12'd2263: chroma9 = 9'b010000110;
        12'd2264: chroma9 = 9'b010001000;
        12'd2265: chroma9 = 9'b010001010;
        12'd2266: chroma9 = 9'b010001100;
        12'd2267: chroma9 = 9'b010001110;
        12'd2268: chroma9 = 9'b010010000;
        12'd2269: chroma9 = 9'b010010011;
        12'd2270: chroma9 = 9'b010010101;
        12'd2271: chroma9 = 9'b010010111;
        12'd2272: chroma9 = 9'b010011010;
        12'd2273: chroma9 = 9'b010011101;
        12'd2274: chroma9 = 9'b010011111;
        12'd2275: chroma9 = 9'b010100010;
        12'd2276: chroma9 = 9'b010100101;
        12'd2277: chroma9 = 9'b010100111;
        12'd2278: chroma9 = 9'b010101010;
        12'd2279: chroma9 = 9'b010101101;
        12'd2280: chroma9 = 9'b010110000;
        12'd2281: chroma9 = 9'b010110011;
        12'd2282: chroma9 = 9'b010110110;
        12'd2283: chroma9 = 9'b010111001;
        12'd2284: chroma9 = 9'b010111100;
        12'd2285: chroma9 = 9'b010111111;
        12'd2286: chroma9 = 9'b011000011;
        12'd2287: chroma9 = 9'b011000110;
        12'd2288: chroma9 = 9'b011001001;
        12'd2289: chroma9 = 9'b011001100;
        12'd2290: chroma9 = 9'b011010000;
        12'd2291: chroma9 = 9'b011010011;
        12'd2292: chroma9 = 9'b011010110;
        12'd2293: chroma9 = 9'b011011010;
        12'd2294: chroma9 = 9'b011011101;
        12'd2295: chroma9 = 9'b011100001;
        12'd2296: chroma9 = 9'b011100100;
        12'd2297: chroma9 = 9'b011101000;
        12'd2298: chroma9 = 9'b011101011;
        12'd2299: chroma9 = 9'b011101111;
        12'd2300: chroma9 = 9'b011110010;
        12'd2301: chroma9 = 9'b011110110;
        12'd2302: chroma9 = 9'b011111001;
        12'd2303: chroma9 = 9'b011111101;
        12'd2304: chroma9 = 9'b100000000;
        12'd2305: chroma9 = 9'b100000011;
        12'd2306: chroma9 = 9'b100000111;
        12'd2307: chroma9 = 9'b100001011;
        12'd2308: chroma9 = 9'b100001111;
        12'd2309: chroma9 = 9'b100010011;
        12'd2310: chroma9 = 9'b100010111;
        12'd2311: chroma9 = 9'b100011011;
        12'd2312: chroma9 = 9'b100011111;
        12'd2313: chroma9 = 9'b100100011;
        12'd2314: chroma9 = 9'b100100110;
        12'd2315: chroma9 = 9'b100101010;
        12'd2316: chroma9 = 9'b100101110;
        12'd2317: chroma9 = 9'b100110010;
        12'd2318: chroma9 = 9'b100110101;
        12'd2319: chroma9 = 9'b100111001;
        12'd2320: chroma9 = 9'b100111101;
        12'd2321: chroma9 = 9'b101000000;
        12'd2322: chroma9 = 9'b101000100;
        12'd2323: chroma9 = 9'b101000111;
        12'd2324: chroma9 = 9'b101001011;
        12'd2325: chroma9 = 9'b101001110;
        12'd2326: chroma9 = 9'b101010010;
        12'd2327: chroma9 = 9'b101010101;
        12'd2328: chroma9 = 9'b101011000;
        12'd2329: chroma9 = 9'b101011100;
        12'd2330: chroma9 = 9'b101011111;
        12'd2331: chroma9 = 9'b101100010;
        12'd2332: chroma9 = 9'b101100101;
        12'd2333: chroma9 = 9'b101101000;
        12'd2334: chroma9 = 9'b101101011;
        12'd2335: chroma9 = 9'b101101110;
        12'd2336: chroma9 = 9'b101110001;
        12'd2337: chroma9 = 9'b101110011;
        12'd2338: chroma9 = 9'b101110110;
        12'd2339: chroma9 = 9'b101111001;
        12'd2340: chroma9 = 9'b101111011;
        12'd2341: chroma9 = 9'b101111110;
        12'd2342: chroma9 = 9'b110000000;
        12'd2343: chroma9 = 9'b110000010;
        12'd2344: chroma9 = 9'b110000101;
        12'd2345: chroma9 = 9'b110000111;
        12'd2346: chroma9 = 9'b110001001;
        12'd2347: chroma9 = 9'b110001011;
        12'd2348: chroma9 = 9'b110001101;
        12'd2349: chroma9 = 9'b110001110;
        12'd2350: chroma9 = 9'b110010000;
        12'd2351: chroma9 = 9'b110010010;
        12'd2352: chroma9 = 9'b110010011;
        12'd2353: chroma9 = 9'b110010101;
        12'd2354: chroma9 = 9'b110010110;
        12'd2355: chroma9 = 9'b110010111;
        12'd2356: chroma9 = 9'b110011001;
        12'd2357: chroma9 = 9'b110011010;
        12'd2358: chroma9 = 9'b110011011;
        12'd2359: chroma9 = 9'b110011100;
        12'd2360: chroma9 = 9'b110011100;
        12'd2361: chroma9 = 9'b110011101;
        12'd2362: chroma9 = 9'b110011110;
        12'd2363: chroma9 = 9'b110011110;
        12'd2364: chroma9 = 9'b110011111;
        12'd2365: chroma9 = 9'b110011111;
        12'd2366: chroma9 = 9'b110011111;
        12'd2367: chroma9 = 9'b110011111;
        12'd2368: chroma9 = 9'b110011111;
        12'd2369: chroma9 = 9'b110011111;
        12'd2370: chroma9 = 9'b110011111;
        12'd2371: chroma9 = 9'b110011111;
        12'd2372: chroma9 = 9'b110011111;
        12'd2373: chroma9 = 9'b110011110;
        12'd2374: chroma9 = 9'b110011110;
        12'd2375: chroma9 = 9'b110011101;
        12'd2376: chroma9 = 9'b110011100;
        12'd2377: chroma9 = 9'b110011100;
        12'd2378: chroma9 = 9'b110011011;
        12'd2379: chroma9 = 9'b110011010;
        12'd2380: chroma9 = 9'b110011001;
        12'd2381: chroma9 = 9'b110010111;
        12'd2382: chroma9 = 9'b110010110;
        12'd2383: chroma9 = 9'b110010101;
        12'd2384: chroma9 = 9'b110010011;
        12'd2385: chroma9 = 9'b110010010;
        12'd2386: chroma9 = 9'b110010000;
        12'd2387: chroma9 = 9'b110001110;
        12'd2388: chroma9 = 9'b110001101;
        12'd2389: chroma9 = 9'b110001011;
        12'd2390: chroma9 = 9'b110001001;
        12'd2391: chroma9 = 9'b110000111;
        12'd2392: chroma9 = 9'b110000101;
        12'd2393: chroma9 = 9'b110000010;
        12'd2394: chroma9 = 9'b110000000;
        12'd2395: chroma9 = 9'b101111110;
        12'd2396: chroma9 = 9'b101111011;
        12'd2397: chroma9 = 9'b101111001;
        12'd2398: chroma9 = 9'b101110110;
        12'd2399: chroma9 = 9'b101110011;
        12'd2400: chroma9 = 9'b101110001;
        12'd2401: chroma9 = 9'b101101110;
        12'd2402: chroma9 = 9'b101101011;
        12'd2403: chroma9 = 9'b101101000;
        12'd2404: chroma9 = 9'b101100101;
        12'd2405: chroma9 = 9'b101100010;
        12'd2406: chroma9 = 9'b101011111;
        12'd2407: chroma9 = 9'b101011100;
        12'd2408: chroma9 = 9'b101011000;
        12'd2409: chroma9 = 9'b101010101;
        12'd2410: chroma9 = 9'b101010010;
        12'd2411: chroma9 = 9'b101001110;
        12'd2412: chroma9 = 9'b101001011;
        12'd2413: chroma9 = 9'b101000111;
        12'd2414: chroma9 = 9'b101000100;
        12'd2415: chroma9 = 9'b101000000;
        12'd2416: chroma9 = 9'b100111101;
        12'd2417: chroma9 = 9'b100111001;
        12'd2418: chroma9 = 9'b100110101;
        12'd2419: chroma9 = 9'b100110010;
        12'd2420: chroma9 = 9'b100101110;
        12'd2421: chroma9 = 9'b100101010;
        12'd2422: chroma9 = 9'b100100110;
        12'd2423: chroma9 = 9'b100100011;
        12'd2424: chroma9 = 9'b100011111;
        12'd2425: chroma9 = 9'b100011011;
        12'd2426: chroma9 = 9'b100010111;
        12'd2427: chroma9 = 9'b100010011;
        12'd2428: chroma9 = 9'b100001111;
        12'd2429: chroma9 = 9'b100001011;
        12'd2430: chroma9 = 9'b100000111;
        12'd2431: chroma9 = 9'b100000011;
        12'd2432: chroma9 = 9'b100000000;
        12'd2433: chroma9 = 9'b011111101;
        12'd2434: chroma9 = 9'b011111001;
        12'd2435: chroma9 = 9'b011110101;
        12'd2436: chroma9 = 9'b011110001;
        12'd2437: chroma9 = 9'b011101101;
        12'd2438: chroma9 = 9'b011101001;
        12'd2439: chroma9 = 9'b011100101;
        12'd2440: chroma9 = 9'b011100001;
        12'd2441: chroma9 = 9'b011011101;
        12'd2442: chroma9 = 9'b011011010;
        12'd2443: chroma9 = 9'b011010110;
        12'd2444: chroma9 = 9'b011010010;
        12'd2445: chroma9 = 9'b011001110;
        12'd2446: chroma9 = 9'b011001011;
        12'd2447: chroma9 = 9'b011000111;
        12'd2448: chroma9 = 9'b011000011;
        12'd2449: chroma9 = 9'b011000000;
        12'd2450: chroma9 = 9'b010111100;
        12'd2451: chroma9 = 9'b010111001;
        12'd2452: chroma9 = 9'b010110101;
        12'd2453: chroma9 = 9'b010110010;
        12'd2454: chroma9 = 9'b010101110;
        12'd2455: chroma9 = 9'b010101011;
        12'd2456: chroma9 = 9'b010101000;
        12'd2457: chroma9 = 9'b010100100;
        12'd2458: chroma9 = 9'b010100001;
        12'd2459: chroma9 = 9'b010011110;
        12'd2460: chroma9 = 9'b010011011;
        12'd2461: chroma9 = 9'b010011000;
        12'd2462: chroma9 = 9'b010010101;
        12'd2463: chroma9 = 9'b010010010;
        12'd2464: chroma9 = 9'b010001111;
        12'd2465: chroma9 = 9'b010001101;
        12'd2466: chroma9 = 9'b010001010;
        12'd2467: chroma9 = 9'b010000111;
        12'd2468: chroma9 = 9'b010000101;
        12'd2469: chroma9 = 9'b010000010;
        12'd2470: chroma9 = 9'b010000000;
        12'd2471: chroma9 = 9'b001111110;
        12'd2472: chroma9 = 9'b001111011;
        12'd2473: chroma9 = 9'b001111001;
        12'd2474: chroma9 = 9'b001110111;
        12'd2475: chroma9 = 9'b001110101;
        12'd2476: chroma9 = 9'b001110011;
        12'd2477: chroma9 = 9'b001110010;
        12'd2478: chroma9 = 9'b001110000;
        12'd2479: chroma9 = 9'b001101110;
        12'd2480: chroma9 = 9'b001101101;
        12'd2481: chroma9 = 9'b001101011;
        12'd2482: chroma9 = 9'b001101010;
        12'd2483: chroma9 = 9'b001101001;
        12'd2484: chroma9 = 9'b001100111;
        12'd2485: chroma9 = 9'b001100110;
        12'd2486: chroma9 = 9'b001100101;
        12'd2487: chroma9 = 9'b001100100;
        12'd2488: chroma9 = 9'b001100100;
        12'd2489: chroma9 = 9'b001100011;
        12'd2490: chroma9 = 9'b001100010;
        12'd2491: chroma9 = 9'b001100010;
        12'd2492: chroma9 = 9'b001100001;
        12'd2493: chroma9 = 9'b001100001;
        12'd2494: chroma9 = 9'b001100001;
        12'd2495: chroma9 = 9'b001100001;
        12'd2496: chroma9 = 9'b001100001;
        12'd2497: chroma9 = 9'b001100001;
        12'd2498: chroma9 = 9'b001100001;
        12'd2499: chroma9 = 9'b001100001;
        12'd2500: chroma9 = 9'b001100001;
        12'd2501: chroma9 = 9'b001100010;
        12'd2502: chroma9 = 9'b001100010;
        12'd2503: chroma9 = 9'b001100011;
        12'd2504: chroma9 = 9'b001100100;
        12'd2505: chroma9 = 9'b001100100;
        12'd2506: chroma9 = 9'b001100101;
        12'd2507: chroma9 = 9'b001100110;
        12'd2508: chroma9 = 9'b001100111;
        12'd2509: chroma9 = 9'b001101001;
        12'd2510: chroma9 = 9'b001101010;
        12'd2511: chroma9 = 9'b001101011;
        12'd2512: chroma9 = 9'b001101101;
        12'd2513: chroma9 = 9'b001101110;
        12'd2514: chroma9 = 9'b001110000;
        12'd2515: chroma9 = 9'b001110010;
        12'd2516: chroma9 = 9'b001110011;
        12'd2517: chroma9 = 9'b001110101;
        12'd2518: chroma9 = 9'b001110111;
        12'd2519: chroma9 = 9'b001111001;
        12'd2520: chroma9 = 9'b001111011;
        12'd2521: chroma9 = 9'b001111110;
        12'd2522: chroma9 = 9'b010000000;
        12'd2523: chroma9 = 9'b010000010;
        12'd2524: chroma9 = 9'b010000101;
        12'd2525: chroma9 = 9'b010000111;
        12'd2526: chroma9 = 9'b010001010;
        12'd2527: chroma9 = 9'b010001101;
        12'd2528: chroma9 = 9'b010001111;
        12'd2529: chroma9 = 9'b010010010;
        12'd2530: chroma9 = 9'b010010101;
        12'd2531: chroma9 = 9'b010011000;
        12'd2532: chroma9 = 9'b010011011;
        12'd2533: chroma9 = 9'b010011110;
        12'd2534: chroma9 = 9'b010100001;
        12'd2535: chroma9 = 9'b010100100;
        12'd2536: chroma9 = 9'b010101000;
        12'd2537: chroma9 = 9'b010101011;
        12'd2538: chroma9 = 9'b010101110;
        12'd2539: chroma9 = 9'b010110010;
        12'd2540: chroma9 = 9'b010110101;
        12'd2541: chroma9 = 9'b010111001;
        12'd2542: chroma9 = 9'b010111100;
        12'd2543: chroma9 = 9'b011000000;
        12'd2544: chroma9 = 9'b011000011;
        12'd2545: chroma9 = 9'b011000111;
        12'd2546: chroma9 = 9'b011001011;
        12'd2547: chroma9 = 9'b011001110;
        12'd2548: chroma9 = 9'b011010010;
        12'd2549: chroma9 = 9'b011010110;
        12'd2550: chroma9 = 9'b011011010;
        12'd2551: chroma9 = 9'b011011101;
        12'd2552: chroma9 = 9'b011100001;
        12'd2553: chroma9 = 9'b011100101;
        12'd2554: chroma9 = 9'b011101001;
        12'd2555: chroma9 = 9'b011101101;
        12'd2556: chroma9 = 9'b011110001;
        12'd2557: chroma9 = 9'b011110101;
        12'd2558: chroma9 = 9'b011111001;
        12'd2559: chroma9 = 9'b011111101;
        12'd2560: chroma9 = 9'b100000000;
        12'd2561: chroma9 = 9'b100000100;
        12'd2562: chroma9 = 9'b100001000;
        12'd2563: chroma9 = 9'b100001100;
        12'd2564: chroma9 = 9'b100010001;
        12'd2565: chroma9 = 9'b100010101;
        12'd2566: chroma9 = 9'b100011001;
        12'd2567: chroma9 = 9'b100011101;
        12'd2568: chroma9 = 9'b100100010;
        12'd2569: chroma9 = 9'b100100110;
        12'd2570: chroma9 = 9'b100101010;
        12'd2571: chroma9 = 9'b100101110;
        12'd2572: chroma9 = 9'b100110010;
        12'd2573: chroma9 = 9'b100110110;
        12'd2574: chroma9 = 9'b100111010;
        12'd2575: chroma9 = 9'b100111110;
        12'd2576: chroma9 = 9'b101000010;
        12'd2577: chroma9 = 9'b101000110;
        12'd2578: chroma9 = 9'b101001010;
        12'd2579: chroma9 = 9'b101001110;
        12'd2580: chroma9 = 9'b101010010;
        12'd2581: chroma9 = 9'b101010110;
        12'd2582: chroma9 = 9'b101011001;
        12'd2583: chroma9 = 9'b101011101;
        12'd2584: chroma9 = 9'b101100001;
        12'd2585: chroma9 = 9'b101100100;
        12'd2586: chroma9 = 9'b101101000;
        12'd2587: chroma9 = 9'b101101011;
        12'd2588: chroma9 = 9'b101101111;
        12'd2589: chroma9 = 9'b101110010;
        12'd2590: chroma9 = 9'b101110101;
        12'd2591: chroma9 = 9'b101111000;
        12'd2592: chroma9 = 9'b101111011;
        12'd2593: chroma9 = 9'b101111110;
        12'd2594: chroma9 = 9'b110000001;
        12'd2595: chroma9 = 9'b110000100;
        12'd2596: chroma9 = 9'b110000111;
        12'd2597: chroma9 = 9'b110001001;
        12'd2598: chroma9 = 9'b110001100;
        12'd2599: chroma9 = 9'b110001111;
        12'd2600: chroma9 = 9'b110010001;
        12'd2601: chroma9 = 9'b110010011;
        12'd2602: chroma9 = 9'b110010110;
        12'd2603: chroma9 = 9'b110011000;
        12'd2604: chroma9 = 9'b110011010;
        12'd2605: chroma9 = 9'b110011100;
        12'd2606: chroma9 = 9'b110011110;
        12'd2607: chroma9 = 9'b110011111;
        12'd2608: chroma9 = 9'b110100001;
        12'd2609: chroma9 = 9'b110100011;
        12'd2610: chroma9 = 9'b110100100;
        12'd2611: chroma9 = 9'b110100110;
        12'd2612: chroma9 = 9'b110100111;
        12'd2613: chroma9 = 9'b110101000;
        12'd2614: chroma9 = 9'b110101001;
        12'd2615: chroma9 = 9'b110101010;
        12'd2616: chroma9 = 9'b110101011;
        12'd2617: chroma9 = 9'b110101100;
        12'd2618: chroma9 = 9'b110101101;
        12'd2619: chroma9 = 9'b110101101;
        12'd2620: chroma9 = 9'b110101110;
        12'd2621: chroma9 = 9'b110101110;
        12'd2622: chroma9 = 9'b110101110;
        12'd2623: chroma9 = 9'b110101110;
        12'd2624: chroma9 = 9'b110101110;
        12'd2625: chroma9 = 9'b110101110;
        12'd2626: chroma9 = 9'b110101110;
        12'd2627: chroma9 = 9'b110101110;
        12'd2628: chroma9 = 9'b110101110;
        12'd2629: chroma9 = 9'b110101101;
        12'd2630: chroma9 = 9'b110101101;
        12'd2631: chroma9 = 9'b110101100;
        12'd2632: chroma9 = 9'b110101011;
        12'd2633: chroma9 = 9'b110101010;
        12'd2634: chroma9 = 9'b110101001;
        12'd2635: chroma9 = 9'b110101000;
        12'd2636: chroma9 = 9'b110100111;
        12'd2637: chroma9 = 9'b110100110;
        12'd2638: chroma9 = 9'b110100100;
        12'd2639: chroma9 = 9'b110100011;
        12'd2640: chroma9 = 9'b110100001;
        12'd2641: chroma9 = 9'b110011111;
        12'd2642: chroma9 = 9'b110011110;
        12'd2643: chroma9 = 9'b110011100;
        12'd2644: chroma9 = 9'b110011010;
        12'd2645: chroma9 = 9'b110011000;
        12'd2646: chroma9 = 9'b110010110;
        12'd2647: chroma9 = 9'b110010011;
        12'd2648: chroma9 = 9'b110010001;
        12'd2649: chroma9 = 9'b110001111;
        12'd2650: chroma9 = 9'b110001100;
        12'd2651: chroma9 = 9'b110001001;
        12'd2652: chroma9 = 9'b110000111;
        12'd2653: chroma9 = 9'b110000100;
        12'd2654: chroma9 = 9'b110000001;
        12'd2655: chroma9 = 9'b101111110;
        12'd2656: chroma9 = 9'b101111011;
        12'd2657: chroma9 = 9'b101111000;
        12'd2658: chroma9 = 9'b101110101;
        12'd2659: chroma9 = 9'b101110010;
        12'd2660: chroma9 = 9'b101101111;
        12'd2661: chroma9 = 9'b101101011;
        12'd2662: chroma9 = 9'b101101000;
        12'd2663: chroma9 = 9'b101100100;
        12'd2664: chroma9 = 9'b101100001;
        12'd2665: chroma9 = 9'b101011101;
        12'd2666: chroma9 = 9'b101011001;
        12'd2667: chroma9 = 9'b101010110;
        12'd2668: chroma9 = 9'b101010010;
        12'd2669: chroma9 = 9'b101001110;
        12'd2670: chroma9 = 9'b101001010;
        12'd2671: chroma9 = 9'b101000110;
        12'd2672: chroma9 = 9'b101000010;
        12'd2673: chroma9 = 9'b100111110;
        12'd2674: chroma9 = 9'b100111010;
        12'd2675: chroma9 = 9'b100110110;
        12'd2676: chroma9 = 9'b100110010;
        12'd2677: chroma9 = 9'b100101110;
        12'd2678: chroma9 = 9'b100101010;
        12'd2679: chroma9 = 9'b100100110;
        12'd2680: chroma9 = 9'b100100010;
        12'd2681: chroma9 = 9'b100011101;
        12'd2682: chroma9 = 9'b100011001;
        12'd2683: chroma9 = 9'b100010101;
        12'd2684: chroma9 = 9'b100010001;
        12'd2685: chroma9 = 9'b100001100;
        12'd2686: chroma9 = 9'b100001000;
        12'd2687: chroma9 = 9'b100000100;
        12'd2688: chroma9 = 9'b100000000;
        12'd2689: chroma9 = 9'b011111100;
        12'd2690: chroma9 = 9'b011111000;
        12'd2691: chroma9 = 9'b011110100;
        12'd2692: chroma9 = 9'b011101111;
        12'd2693: chroma9 = 9'b011101011;
        12'd2694: chroma9 = 9'b011100111;
        12'd2695: chroma9 = 9'b011100011;
        12'd2696: chroma9 = 9'b011011110;
        12'd2697: chroma9 = 9'b011011010;
        12'd2698: chroma9 = 9'b011010110;
        12'd2699: chroma9 = 9'b011010010;
        12'd2700: chroma9 = 9'b011001110;
        12'd2701: chroma9 = 9'b011001010;
        12'd2702: chroma9 = 9'b011000110;
        12'd2703: chroma9 = 9'b011000010;
        12'd2704: chroma9 = 9'b010111110;
        12'd2705: chroma9 = 9'b010111010;
        12'd2706: chroma9 = 9'b010110110;
        12'd2707: chroma9 = 9'b010110010;
        12'd2708: chroma9 = 9'b010101110;
        12'd2709: chroma9 = 9'b010101010;
        12'd2710: chroma9 = 9'b010100111;
        12'd2711: chroma9 = 9'b010100011;
        12'd2712: chroma9 = 9'b010011111;
        12'd2713: chroma9 = 9'b010011100;
        12'd2714: chroma9 = 9'b010011000;
        12'd2715: chroma9 = 9'b010010101;
        12'd2716: chroma9 = 9'b010010001;
        12'd2717: chroma9 = 9'b010001110;
        12'd2718: chroma9 = 9'b010001011;
        12'd2719: chroma9 = 9'b010001000;
        12'd2720: chroma9 = 9'b010000101;
        12'd2721: chroma9 = 9'b010000010;
        12'd2722: chroma9 = 9'b001111111;
        12'd2723: chroma9 = 9'b001111100;
        12'd2724: chroma9 = 9'b001111001;
        12'd2725: chroma9 = 9'b001110111;
        12'd2726: chroma9 = 9'b001110100;
        12'd2727: chroma9 = 9'b001110001;
        12'd2728: chroma9 = 9'b001101111;
        12'd2729: chroma9 = 9'b001101101;
        12'd2730: chroma9 = 9'b001101010;
        12'd2731: chroma9 = 9'b001101000;
        12'd2732: chroma9 = 9'b001100110;
        12'd2733: chroma9 = 9'b001100100;
        12'd2734: chroma9 = 9'b001100010;
        12'd2735: chroma9 = 9'b001100001;
        12'd2736: chroma9 = 9'b001011111;
        12'd2737: chroma9 = 9'b001011101;
        12'd2738: chroma9 = 9'b001011100;
        12'd2739: chroma9 = 9'b001011010;
        12'd2740: chroma9 = 9'b001011001;
        12'd2741: chroma9 = 9'b001011000;
        12'd2742: chroma9 = 9'b001010111;
        12'd2743: chroma9 = 9'b001010110;
        12'd2744: chroma9 = 9'b001010101;
        12'd2745: chroma9 = 9'b001010100;
        12'd2746: chroma9 = 9'b001010011;
        12'd2747: chroma9 = 9'b001010011;
        12'd2748: chroma9 = 9'b001010010;
        12'd2749: chroma9 = 9'b001010010;
        12'd2750: chroma9 = 9'b001010010;
        12'd2751: chroma9 = 9'b001010010;
        12'd2752: chroma9 = 9'b001010010;
        12'd2753: chroma9 = 9'b001010010;
        12'd2754: chroma9 = 9'b001010010;
        12'd2755: chroma9 = 9'b001010010;
        12'd2756: chroma9 = 9'b001010010;
        12'd2757: chroma9 = 9'b001010011;
        12'd2758: chroma9 = 9'b001010011;
        12'd2759: chroma9 = 9'b001010100;
        12'd2760: chroma9 = 9'b001010101;
        12'd2761: chroma9 = 9'b001010110;
        12'd2762: chroma9 = 9'b001010111;
        12'd2763: chroma9 = 9'b001011000;
        12'd2764: chroma9 = 9'b001011001;
        12'd2765: chroma9 = 9'b001011010;
        12'd2766: chroma9 = 9'b001011100;
        12'd2767: chroma9 = 9'b001011101;
        12'd2768: chroma9 = 9'b001011111;
        12'd2769: chroma9 = 9'b001100001;
        12'd2770: chroma9 = 9'b001100010;
        12'd2771: chroma9 = 9'b001100100;
        12'd2772: chroma9 = 9'b001100110;
        12'd2773: chroma9 = 9'b001101000;
        12'd2774: chroma9 = 9'b001101010;
        12'd2775: chroma9 = 9'b001101101;
        12'd2776: chroma9 = 9'b001101111;
        12'd2777: chroma9 = 9'b001110001;
        12'd2778: chroma9 = 9'b001110100;
        12'd2779: chroma9 = 9'b001110111;
        12'd2780: chroma9 = 9'b001111001;
        12'd2781: chroma9 = 9'b001111100;
        12'd2782: chroma9 = 9'b001111111;
        12'd2783: chroma9 = 9'b010000010;
        12'd2784: chroma9 = 9'b010000101;
        12'd2785: chroma9 = 9'b010001000;
        12'd2786: chroma9 = 9'b010001011;
        12'd2787: chroma9 = 9'b010001110;
        12'd2788: chroma9 = 9'b010010001;
        12'd2789: chroma9 = 9'b010010101;
        12'd2790: chroma9 = 9'b010011000;
        12'd2791: chroma9 = 9'b010011100;
        12'd2792: chroma9 = 9'b010011111;
        12'd2793: chroma9 = 9'b010100011;
        12'd2794: chroma9 = 9'b010100111;
        12'd2795: chroma9 = 9'b010101010;
        12'd2796: chroma9 = 9'b010101110;
        12'd2797: chroma9 = 9'b010110010;
        12'd2798: chroma9 = 9'b010110110;
        12'd2799: chroma9 = 9'b010111010;
        12'd2800: chroma9 = 9'b010111110;
        12'd2801: chroma9 = 9'b011000010;
        12'd2802: chroma9 = 9'b011000110;
        12'd2803: chroma9 = 9'b011001010;
        12'd2804: chroma9 = 9'b011001110;
        12'd2805: chroma9 = 9'b011010010;
        12'd2806: chroma9 = 9'b011010110;
        12'd2807: chroma9 = 9'b011011010;
        12'd2808: chroma9 = 9'b011011110;
        12'd2809: chroma9 = 9'b011100011;
        12'd2810: chroma9 = 9'b011100111;
        12'd2811: chroma9 = 9'b011101011;
        12'd2812: chroma9 = 9'b011101111;
        12'd2813: chroma9 = 9'b011110100;
        12'd2814: chroma9 = 9'b011111000;
        12'd2815: chroma9 = 9'b011111100;
        12'd2816: chroma9 = 9'b100000000;
        12'd2817: chroma9 = 9'b100000100;
        12'd2818: chroma9 = 9'b100001001;
        12'd2819: chroma9 = 9'b100001101;
        12'd2820: chroma9 = 9'b100010010;
        12'd2821: chroma9 = 9'b100010111;
        12'd2822: chroma9 = 9'b100011011;
        12'd2823: chroma9 = 9'b100100000;
        12'd2824: chroma9 = 9'b100100101;
        12'd2825: chroma9 = 9'b100101001;
        12'd2826: chroma9 = 9'b100101110;
        12'd2827: chroma9 = 9'b100110010;
        12'd2828: chroma9 = 9'b100110111;
        12'd2829: chroma9 = 9'b100111011;
        12'd2830: chroma9 = 9'b101000000;
        12'd2831: chroma9 = 9'b101000100;
        12'd2832: chroma9 = 9'b101001000;
        12'd2833: chroma9 = 9'b101001100;
        12'd2834: chroma9 = 9'b101010001;
        12'd2835: chroma9 = 9'b101010101;
        12'd2836: chroma9 = 9'b101011001;
        12'd2837: chroma9 = 9'b101011101;
        12'd2838: chroma9 = 9'b101100001;
        12'd2839: chroma9 = 9'b101100101;
        12'd2840: chroma9 = 9'b101101001;
        12'd2841: chroma9 = 9'b101101101;
        12'd2842: chroma9 = 9'b101110001;
        12'd2843: chroma9 = 9'b101110100;
        12'd2844: chroma9 = 9'b101111000;
        12'd2845: chroma9 = 9'b101111100;
        12'd2846: chroma9 = 9'b101111111;
        12'd2847: chroma9 = 9'b110000011;
        12'd2848: chroma9 = 9'b110000110;
        12'd2849: chroma9 = 9'b110001001;
        12'd2850: chroma9 = 9'b110001100;
        12'd2851: chroma9 = 9'b110001111;
        12'd2852: chroma9 = 9'b110010010;
        12'd2853: chroma9 = 9'b110010101;
        12'd2854: chroma9 = 9'b110011000;
        12'd2855: chroma9 = 9'b110011011;
        12'd2856: chroma9 = 9'b110011101;
        12'd2857: chroma9 = 9'b110100000;
        12'd2858: chroma9 = 9'b110100010;
        12'd2859: chroma9 = 9'b110100101;
        12'd2860: chroma9 = 9'b110100111;
        12'd2861: chroma9 = 9'b110101001;
        12'd2862: chroma9 = 9'b110101011;
        12'd2863: chroma9 = 9'b110101101;
        12'd2864: chroma9 = 9'b110101111;
        12'd2865: chroma9 = 9'b110110001;
        12'd2866: chroma9 = 9'b110110010;
        12'd2867: chroma9 = 9'b110110100;
        12'd2868: chroma9 = 9'b110110101;
        12'd2869: chroma9 = 9'b110110111;
        12'd2870: chroma9 = 9'b110111000;
        12'd2871: chroma9 = 9'b110111001;
        12'd2872: chroma9 = 9'b110111010;
        12'd2873: chroma9 = 9'b110111011;
        12'd2874: chroma9 = 9'b110111011;
        12'd2875: chroma9 = 9'b110111100;
        12'd2876: chroma9 = 9'b110111101;
        12'd2877: chroma9 = 9'b110111101;
        12'd2878: chroma9 = 9'b110111101;
        12'd2879: chroma9 = 9'b110111101;
        12'd2880: chroma9 = 9'b110111101;
        12'd2881: chroma9 = 9'b110111101;
        12'd2882: chroma9 = 9'b110111101;
        12'd2883: chroma9 = 9'b110111101;
        12'd2884: chroma9 = 9'b110111101;
        12'd2885: chroma9 = 9'b110111100;
        12'd2886: chroma9 = 9'b110111011;
        12'd2887: chroma9 = 9'b110111011;
        12'd2888: chroma9 = 9'b110111010;
        12'd2889: chroma9 = 9'b110111001;
        12'd2890: chroma9 = 9'b110111000;
        12'd2891: chroma9 = 9'b110110111;
        12'd2892: chroma9 = 9'b110110101;
        12'd2893: chroma9 = 9'b110110100;
        12'd2894: chroma9 = 9'b110110010;
        12'd2895: chroma9 = 9'b110110001;
        12'd2896: chroma9 = 9'b110101111;
        12'd2897: chroma9 = 9'b110101101;
        12'd2898: chroma9 = 9'b110101011;
        12'd2899: chroma9 = 9'b110101001;
        12'd2900: chroma9 = 9'b110100111;
        12'd2901: chroma9 = 9'b110100101;
        12'd2902: chroma9 = 9'b110100010;
        12'd2903: chroma9 = 9'b110100000;
        12'd2904: chroma9 = 9'b110011101;
        12'd2905: chroma9 = 9'b110011011;
        12'd2906: chroma9 = 9'b110011000;
        12'd2907: chroma9 = 9'b110010101;
        12'd2908: chroma9 = 9'b110010010;
        12'd2909: chroma9 = 9'b110001111;
        12'd2910: chroma9 = 9'b110001100;
        12'd2911: chroma9 = 9'b110001001;
        12'd2912: chroma9 = 9'b110000110;
        12'd2913: chroma9 = 9'b110000011;
        12'd2914: chroma9 = 9'b101111111;
        12'd2915: chroma9 = 9'b101111100;
        12'd2916: chroma9 = 9'b101111000;
        12'd2917: chroma9 = 9'b101110100;
        12'd2918: chroma9 = 9'b101110001;
        12'd2919: chroma9 = 9'b101101101;
        12'd2920: chroma9 = 9'b101101001;
        12'd2921: chroma9 = 9'b101100101;
        12'd2922: chroma9 = 9'b101100001;
        12'd2923: chroma9 = 9'b101011101;
        12'd2924: chroma9 = 9'b101011001;
        12'd2925: chroma9 = 9'b101010101;
        12'd2926: chroma9 = 9'b101010001;
        12'd2927: chroma9 = 9'b101001100;
        12'd2928: chroma9 = 9'b101001000;
        12'd2929: chroma9 = 9'b101000100;
        12'd2930: chroma9 = 9'b101000000;
        12'd2931: chroma9 = 9'b100111011;
        12'd2932: chroma9 = 9'b100110111;
        12'd2933: chroma9 = 9'b100110010;
        12'd2934: chroma9 = 9'b100101110;
        12'd2935: chroma9 = 9'b100101001;
        12'd2936: chroma9 = 9'b100100101;
        12'd2937: chroma9 = 9'b100100000;
        12'd2938: chroma9 = 9'b100011011;
        12'd2939: chroma9 = 9'b100010111;
        12'd2940: chroma9 = 9'b100010010;
        12'd2941: chroma9 = 9'b100001101;
        12'd2942: chroma9 = 9'b100001001;
        12'd2943: chroma9 = 9'b100000100;
        12'd2944: chroma9 = 9'b100000000;
        12'd2945: chroma9 = 9'b011111100;
        12'd2946: chroma9 = 9'b011110111;
        12'd2947: chroma9 = 9'b011110011;
        12'd2948: chroma9 = 9'b011101110;
        12'd2949: chroma9 = 9'b011101001;
        12'd2950: chroma9 = 9'b011100101;
        12'd2951: chroma9 = 9'b011100000;
        12'd2952: chroma9 = 9'b011011011;
        12'd2953: chroma9 = 9'b011010111;
        12'd2954: chroma9 = 9'b011010010;
        12'd2955: chroma9 = 9'b011001110;
        12'd2956: chroma9 = 9'b011001001;
        12'd2957: chroma9 = 9'b011000101;
        12'd2958: chroma9 = 9'b011000000;
        12'd2959: chroma9 = 9'b010111100;
        12'd2960: chroma9 = 9'b010111000;
        12'd2961: chroma9 = 9'b010110100;
        12'd2962: chroma9 = 9'b010101111;
        12'd2963: chroma9 = 9'b010101011;
        12'd2964: chroma9 = 9'b010100111;
        12'd2965: chroma9 = 9'b010100011;
        12'd2966: chroma9 = 9'b010011111;
        12'd2967: chroma9 = 9'b010011011;
        12'd2968: chroma9 = 9'b010010111;
        12'd2969: chroma9 = 9'b010010011;
        12'd2970: chroma9 = 9'b010001111;
        12'd2971: chroma9 = 9'b010001100;
        12'd2972: chroma9 = 9'b010001000;
        12'd2973: chroma9 = 9'b010000100;
        12'd2974: chroma9 = 9'b010000001;
        12'd2975: chroma9 = 9'b001111101;
        12'd2976: chroma9 = 9'b001111010;
        12'd2977: chroma9 = 9'b001110111;
        12'd2978: chroma9 = 9'b001110100;
        12'd2979: chroma9 = 9'b001110001;
        12'd2980: chroma9 = 9'b001101110;
        12'd2981: chroma9 = 9'b001101011;
        12'd2982: chroma9 = 9'b001101000;
        12'd2983: chroma9 = 9'b001100101;
        12'd2984: chroma9 = 9'b001100011;
        12'd2985: chroma9 = 9'b001100000;
        12'd2986: chroma9 = 9'b001011110;
        12'd2987: chroma9 = 9'b001011011;
        12'd2988: chroma9 = 9'b001011001;
        12'd2989: chroma9 = 9'b001010111;
        12'd2990: chroma9 = 9'b001010101;
        12'd2991: chroma9 = 9'b001010011;
        12'd2992: chroma9 = 9'b001010001;
        12'd2993: chroma9 = 9'b001001111;
        12'd2994: chroma9 = 9'b001001110;
        12'd2995: chroma9 = 9'b001001100;
        12'd2996: chroma9 = 9'b001001011;
        12'd2997: chroma9 = 9'b001001001;
        12'd2998: chroma9 = 9'b001001000;
        12'd2999: chroma9 = 9'b001000111;
        12'd3000: chroma9 = 9'b001000110;
        12'd3001: chroma9 = 9'b001000101;
        12'd3002: chroma9 = 9'b001000101;
        12'd3003: chroma9 = 9'b001000100;
        12'd3004: chroma9 = 9'b001000011;
        12'd3005: chroma9 = 9'b001000011;
        12'd3006: chroma9 = 9'b001000011;
        12'd3007: chroma9 = 9'b001000011;
        12'd3008: chroma9 = 9'b001000011;
        12'd3009: chroma9 = 9'b001000011;
        12'd3010: chroma9 = 9'b001000011;
        12'd3011: chroma9 = 9'b001000011;
        12'd3012: chroma9 = 9'b001000011;
        12'd3013: chroma9 = 9'b001000100;
        12'd3014: chroma9 = 9'b001000101;
        12'd3015: chroma9 = 9'b001000101;
        12'd3016: chroma9 = 9'b001000110;
        12'd3017: chroma9 = 9'b001000111;
        12'd3018: chroma9 = 9'b001001000;
        12'd3019: chroma9 = 9'b001001001;
        12'd3020: chroma9 = 9'b001001011;
        12'd3021: chroma9 = 9'b001001100;
        12'd3022: chroma9 = 9'b001001110;
        12'd3023: chroma9 = 9'b001001111;
        12'd3024: chroma9 = 9'b001010001;
        12'd3025: chroma9 = 9'b001010011;
        12'd3026: chroma9 = 9'b001010101;
        12'd3027: chroma9 = 9'b001010111;
        12'd3028: chroma9 = 9'b001011001;
        12'd3029: chroma9 = 9'b001011011;
        12'd3030: chroma9 = 9'b001011110;
        12'd3031: chroma9 = 9'b001100000;
        12'd3032: chroma9 = 9'b001100011;
        12'd3033: chroma9 = 9'b001100101;
        12'd3034: chroma9 = 9'b001101000;
        12'd3035: chroma9 = 9'b001101011;
        12'd3036: chroma9 = 9'b001101110;
        12'd3037: chroma9 = 9'b001110001;
        12'd3038: chroma9 = 9'b001110100;
        12'd3039: chroma9 = 9'b001110111;
        12'd3040: chroma9 = 9'b001111010;
        12'd3041: chroma9 = 9'b001111101;
        12'd3042: chroma9 = 9'b010000001;
        12'd3043: chroma9 = 9'b010000100;
        12'd3044: chroma9 = 9'b010001000;
        12'd3045: chroma9 = 9'b010001100;
        12'd3046: chroma9 = 9'b010001111;
        12'd3047: chroma9 = 9'b010010011;
        12'd3048: chroma9 = 9'b010010111;
        12'd3049: chroma9 = 9'b010011011;
        12'd3050: chroma9 = 9'b010011111;
        12'd3051: chroma9 = 9'b010100011;
        12'd3052: chroma9 = 9'b010100111;
        12'd3053: chroma9 = 9'b010101011;
        12'd3054: chroma9 = 9'b010101111;
        12'd3055: chroma9 = 9'b010110100;
        12'd3056: chroma9 = 9'b010111000;
        12'd3057: chroma9 = 9'b010111100;
        12'd3058: chroma9 = 9'b011000000;
        12'd3059: chroma9 = 9'b011000101;
        12'd3060: chroma9 = 9'b011001001;
        12'd3061: chroma9 = 9'b011001110;
        12'd3062: chroma9 = 9'b011010010;
        12'd3063: chroma9 = 9'b011010111;
        12'd3064: chroma9 = 9'b011011011;
        12'd3065: chroma9 = 9'b011100000;
        12'd3066: chroma9 = 9'b011100101;
        12'd3067: chroma9 = 9'b011101001;
        12'd3068: chroma9 = 9'b011101110;
        12'd3069: chroma9 = 9'b011110011;
        12'd3070: chroma9 = 9'b011110111;
        12'd3071: chroma9 = 9'b011111100;
        12'd3072: chroma9 = 9'b100000000;
        12'd3073: chroma9 = 9'b100000101;
        12'd3074: chroma9 = 9'b100001010;
        12'd3075: chroma9 = 9'b100001111;
        12'd3076: chroma9 = 9'b100010100;
        12'd3077: chroma9 = 9'b100011001;
        12'd3078: chroma9 = 9'b100011110;
        12'd3079: chroma9 = 9'b100100011;
        12'd3080: chroma9 = 9'b100100111;
        12'd3081: chroma9 = 9'b100101100;
        12'd3082: chroma9 = 9'b100110001;
        12'd3083: chroma9 = 9'b100110110;
        12'd3084: chroma9 = 9'b100111011;
        12'd3085: chroma9 = 9'b101000000;
        12'd3086: chroma9 = 9'b101000101;
        12'd3087: chroma9 = 9'b101001001;
        12'd3088: chroma9 = 9'b101001110;
        12'd3089: chroma9 = 9'b101010011;
        12'd3090: chroma9 = 9'b101010111;
        12'd3091: chroma9 = 9'b101011100;
        12'd3092: chroma9 = 9'b101100000;
        12'd3093: chroma9 = 9'b101100101;
        12'd3094: chroma9 = 9'b101101001;
        12'd3095: chroma9 = 9'b101101101;
        12'd3096: chroma9 = 9'b101110001;
        12'd3097: chroma9 = 9'b101110110;
        12'd3098: chroma9 = 9'b101111010;
        12'd3099: chroma9 = 9'b101111110;
        12'd3100: chroma9 = 9'b110000010;
        12'd3101: chroma9 = 9'b110000101;
        12'd3102: chroma9 = 9'b110001001;
        12'd3103: chroma9 = 9'b110001101;
        12'd3104: chroma9 = 9'b110010000;
        12'd3105: chroma9 = 9'b110010100;
        12'd3106: chroma9 = 9'b110010111;
        12'd3107: chroma9 = 9'b110011011;
        12'd3108: chroma9 = 9'b110011110;
        12'd3109: chroma9 = 9'b110100001;
        12'd3110: chroma9 = 9'b110100100;
        12'd3111: chroma9 = 9'b110100111;
        12'd3112: chroma9 = 9'b110101010;
        12'd3113: chroma9 = 9'b110101101;
        12'd3114: chroma9 = 9'b110101111;
        12'd3115: chroma9 = 9'b110110010;
        12'd3116: chroma9 = 9'b110110100;
        12'd3117: chroma9 = 9'b110110111;
        12'd3118: chroma9 = 9'b110111001;
        12'd3119: chroma9 = 9'b110111011;
        12'd3120: chroma9 = 9'b110111101;
        12'd3121: chroma9 = 9'b110111111;
        12'd3122: chroma9 = 9'b111000001;
        12'd3123: chroma9 = 9'b111000010;
        12'd3124: chroma9 = 9'b111000100;
        12'd3125: chroma9 = 9'b111000101;
        12'd3126: chroma9 = 9'b111000110;
        12'd3127: chroma9 = 9'b111001000;
        12'd3128: chroma9 = 9'b111001001;
        12'd3129: chroma9 = 9'b111001001;
        12'd3130: chroma9 = 9'b111001010;
        12'd3131: chroma9 = 9'b111001011;
        12'd3132: chroma9 = 9'b111001100;
        12'd3133: chroma9 = 9'b111001100;
        12'd3134: chroma9 = 9'b111001100;
        12'd3135: chroma9 = 9'b111001100;
        12'd3136: chroma9 = 9'b111001100;
        12'd3137: chroma9 = 9'b111001100;
        12'd3138: chroma9 = 9'b111001100;
        12'd3139: chroma9 = 9'b111001100;
        12'd3140: chroma9 = 9'b111001100;
        12'd3141: chroma9 = 9'b111001011;
        12'd3142: chroma9 = 9'b111001010;
        12'd3143: chroma9 = 9'b111001001;
        12'd3144: chroma9 = 9'b111001001;
        12'd3145: chroma9 = 9'b111001000;
        12'd3146: chroma9 = 9'b111000110;
        12'd3147: chroma9 = 9'b111000101;
        12'd3148: chroma9 = 9'b111000100;
        12'd3149: chroma9 = 9'b111000010;
        12'd3150: chroma9 = 9'b111000001;
        12'd3151: chroma9 = 9'b110111111;
        12'd3152: chroma9 = 9'b110111101;
        12'd3153: chroma9 = 9'b110111011;
        12'd3154: chroma9 = 9'b110111001;
        12'd3155: chroma9 = 9'b110110111;
        12'd3156: chroma9 = 9'b110110100;
        12'd3157: chroma9 = 9'b110110010;
        12'd3158: chroma9 = 9'b110101111;
        12'd3159: chroma9 = 9'b110101101;
        12'd3160: chroma9 = 9'b110101010;
        12'd3161: chroma9 = 9'b110100111;
        12'd3162: chroma9 = 9'b110100100;
        12'd3163: chroma9 = 9'b110100001;
        12'd3164: chroma9 = 9'b110011110;
        12'd3165: chroma9 = 9'b110011011;
        12'd3166: chroma9 = 9'b110010111;
        12'd3167: chroma9 = 9'b110010100;
        12'd3168: chroma9 = 9'b110010000;
        12'd3169: chroma9 = 9'b110001101;
        12'd3170: chroma9 = 9'b110001001;
        12'd3171: chroma9 = 9'b110000101;
        12'd3172: chroma9 = 9'b110000010;
        12'd3173: chroma9 = 9'b101111110;
        12'd3174: chroma9 = 9'b101111010;
        12'd3175: chroma9 = 9'b101110110;
        12'd3176: chroma9 = 9'b101110001;
        12'd3177: chroma9 = 9'b101101101;
        12'd3178: chroma9 = 9'b101101001;
        12'd3179: chroma9 = 9'b101100101;
        12'd3180: chroma9 = 9'b101100000;
        12'd3181: chroma9 = 9'b101011100;
        12'd3182: chroma9 = 9'b101010111;
        12'd3183: chroma9 = 9'b101010011;
        12'd3184: chroma9 = 9'b101001110;
        12'd3185: chroma9 = 9'b101001001;
        12'd3186: chroma9 = 9'b101000101;
        12'd3187: chroma9 = 9'b101000000;
        12'd3188: chroma9 = 9'b100111011;
        12'd3189: chroma9 = 9'b100110110;
        12'd3190: chroma9 = 9'b100110001;
        12'd3191: chroma9 = 9'b100101100;
        12'd3192: chroma9 = 9'b100100111;
        12'd3193: chroma9 = 9'b100100011;
        12'd3194: chroma9 = 9'b100011110;
        12'd3195: chroma9 = 9'b100011001;
        12'd3196: chroma9 = 9'b100010100;
        12'd3197: chroma9 = 9'b100001111;
        12'd3198: chroma9 = 9'b100001010;
        12'd3199: chroma9 = 9'b100000101;
        12'd3200: chroma9 = 9'b100000000;
        12'd3201: chroma9 = 9'b011111011;
        12'd3202: chroma9 = 9'b011110110;
        12'd3203: chroma9 = 9'b011110001;
        12'd3204: chroma9 = 9'b011101100;
        12'd3205: chroma9 = 9'b011100111;
        12'd3206: chroma9 = 9'b011100010;
        12'd3207: chroma9 = 9'b011011101;
        12'd3208: chroma9 = 9'b011011001;
        12'd3209: chroma9 = 9'b011010100;
        12'd3210: chroma9 = 9'b011001111;
        12'd3211: chroma9 = 9'b011001010;
        12'd3212: chroma9 = 9'b011000101;
        12'd3213: chroma9 = 9'b011000000;
        12'd3214: chroma9 = 9'b010111011;
        12'd3215: chroma9 = 9'b010110111;
        12'd3216: chroma9 = 9'b010110010;
        12'd3217: chroma9 = 9'b010101101;
        12'd3218: chroma9 = 9'b010101001;
        12'd3219: chroma9 = 9'b010100100;
        12'd3220: chroma9 = 9'b010100000;
        12'd3221: chroma9 = 9'b010011011;
        12'd3222: chroma9 = 9'b010010111;
        12'd3223: chroma9 = 9'b010010011;
        12'd3224: chroma9 = 9'b010001111;
        12'd3225: chroma9 = 9'b010001010;
        12'd3226: chroma9 = 9'b010000110;
        12'd3227: chroma9 = 9'b010000010;
        12'd3228: chroma9 = 9'b001111110;
        12'd3229: chroma9 = 9'b001111011;
        12'd3230: chroma9 = 9'b001110111;
        12'd3231: chroma9 = 9'b001110011;
        12'd3232: chroma9 = 9'b001110000;
        12'd3233: chroma9 = 9'b001101100;
        12'd3234: chroma9 = 9'b001101001;
        12'd3235: chroma9 = 9'b001100101;
        12'd3236: chroma9 = 9'b001100010;
        12'd3237: chroma9 = 9'b001011111;
        12'd3238: chroma9 = 9'b001011100;
        12'd3239: chroma9 = 9'b001011001;
        12'd3240: chroma9 = 9'b001010110;
        12'd3241: chroma9 = 9'b001010011;
        12'd3242: chroma9 = 9'b001010001;
        12'd3243: chroma9 = 9'b001001110;
        12'd3244: chroma9 = 9'b001001100;
        12'd3245: chroma9 = 9'b001001001;
        12'd3246: chroma9 = 9'b001000111;
        12'd3247: chroma9 = 9'b001000101;
        12'd3248: chroma9 = 9'b001000011;
        12'd3249: chroma9 = 9'b001000001;
        12'd3250: chroma9 = 9'b000111111;
        12'd3251: chroma9 = 9'b000111110;
        12'd3252: chroma9 = 9'b000111100;
        12'd3253: chroma9 = 9'b000111011;
        12'd3254: chroma9 = 9'b000111010;
        12'd3255: chroma9 = 9'b000111000;
        12'd3256: chroma9 = 9'b000110111;
        12'd3257: chroma9 = 9'b000110111;
        12'd3258: chroma9 = 9'b000110110;
        12'd3259: chroma9 = 9'b000110101;
        12'd3260: chroma9 = 9'b000110100;
        12'd3261: chroma9 = 9'b000110100;
        12'd3262: chroma9 = 9'b000110100;
        12'd3263: chroma9 = 9'b000110100;
        12'd3264: chroma9 = 9'b000110100;
        12'd3265: chroma9 = 9'b000110100;
        12'd3266: chroma9 = 9'b000110100;
        12'd3267: chroma9 = 9'b000110100;
        12'd3268: chroma9 = 9'b000110100;
        12'd3269: chroma9 = 9'b000110101;
        12'd3270: chroma9 = 9'b000110110;
        12'd3271: chroma9 = 9'b000110111;
        12'd3272: chroma9 = 9'b000110111;
        12'd3273: chroma9 = 9'b000111000;
        12'd3274: chroma9 = 9'b000111010;
        12'd3275: chroma9 = 9'b000111011;
        12'd3276: chroma9 = 9'b000111100;
        12'd3277: chroma9 = 9'b000111110;
        12'd3278: chroma9 = 9'b000111111;
        12'd3279: chroma9 = 9'b001000001;
        12'd3280: chroma9 = 9'b001000011;
        12'd3281: chroma9 = 9'b001000101;
        12'd3282: chroma9 = 9'b001000111;
        12'd3283: chroma9 = 9'b001001001;
        12'd3284: chroma9 = 9'b001001100;
        12'd3285: chroma9 = 9'b001001110;
        12'd3286: chroma9 = 9'b001010001;
        12'd3287: chroma9 = 9'b001010011;
        12'd3288: chroma9 = 9'b001010110;
        12'd3289: chroma9 = 9'b001011001;
        12'd3290: chroma9 = 9'b001011100;
        12'd3291: chroma9 = 9'b001011111;
        12'd3292: chroma9 = 9'b001100010;
        12'd3293: chroma9 = 9'b001100101;
        12'd3294: chroma9 = 9'b001101001;
        12'd3295: chroma9 = 9'b001101100;
        12'd3296: chroma9 = 9'b001110000;
        12'd3297: chroma9 = 9'b001110011;
        12'd3298: chroma9 = 9'b001110111;
        12'd3299: chroma9 = 9'b001111011;
        12'd3300: chroma9 = 9'b001111110;
        12'd3301: chroma9 = 9'b010000010;
        12'd3302: chroma9 = 9'b010000110;
        12'd3303: chroma9 = 9'b010001010;
        12'd3304: chroma9 = 9'b010001111;
        12'd3305: chroma9 = 9'b010010011;
        12'd3306: chroma9 = 9'b010010111;
        12'd3307: chroma9 = 9'b010011011;
        12'd3308: chroma9 = 9'b010100000;
        12'd3309: chroma9 = 9'b010100100;
        12'd3310: chroma9 = 9'b010101001;
        12'd3311: chroma9 = 9'b010101101;
        12'd3312: chroma9 = 9'b010110010;
        12'd3313: chroma9 = 9'b010110111;
        12'd3314: chroma9 = 9'b010111011;
        12'd3315: chroma9 = 9'b011000000;
        12'd3316: chroma9 = 9'b011000101;
        12'd3317: chroma9 = 9'b011001010;
        12'd3318: chroma9 = 9'b011001111;
        12'd3319: chroma9 = 9'b011010100;
        12'd3320: chroma9 = 9'b011011001;
        12'd3321: chroma9 = 9'b011011101;
        12'd3322: chroma9 = 9'b011100010;
        12'd3323: chroma9 = 9'b011100111;
        12'd3324: chroma9 = 9'b011101100;
        12'd3325: chroma9 = 9'b011110001;
        12'd3326: chroma9 = 9'b011110110;
        12'd3327: chroma9 = 9'b011111011;
        12'd3328: chroma9 = 9'b100000000;
        12'd3329: chroma9 = 9'b100000101;
        12'd3330: chroma9 = 9'b100001010;
        12'd3331: chroma9 = 9'b100010000;
        12'd3332: chroma9 = 9'b100010101;
        12'd3333: chroma9 = 9'b100011010;
        12'd3334: chroma9 = 9'b100100000;
        12'd3335: chroma9 = 9'b100100101;
        12'd3336: chroma9 = 9'b100101010;
        12'd3337: chroma9 = 9'b100110000;
        12'd3338: chroma9 = 9'b100110101;
        12'd3339: chroma9 = 9'b100111010;
        12'd3340: chroma9 = 9'b100111111;
        12'd3341: chroma9 = 9'b101000101;
        12'd3342: chroma9 = 9'b101001010;
        12'd3343: chroma9 = 9'b101001111;
        12'd3344: chroma9 = 9'b101010100;
        12'd3345: chroma9 = 9'b101011001;
        12'd3346: chroma9 = 9'b101011110;
        12'd3347: chroma9 = 9'b101100010;
        12'd3348: chroma9 = 9'b101100111;
        12'd3349: chroma9 = 9'b101101100;
        12'd3350: chroma9 = 9'b101110001;
        12'd3351: chroma9 = 9'b101110101;
        12'd3352: chroma9 = 9'b101111010;
        12'd3353: chroma9 = 9'b101111110;
        12'd3354: chroma9 = 9'b110000011;
        12'd3355: chroma9 = 9'b110000111;
        12'd3356: chroma9 = 9'b110001011;
        12'd3357: chroma9 = 9'b110001111;
        12'd3358: chroma9 = 9'b110010011;
        12'd3359: chroma9 = 9'b110010111;
        12'd3360: chroma9 = 9'b110011011;
        12'd3361: chroma9 = 9'b110011111;
        12'd3362: chroma9 = 9'b110100011;
        12'd3363: chroma9 = 9'b110100110;
        12'd3364: chroma9 = 9'b110101010;
        12'd3365: chroma9 = 9'b110101101;
        12'd3366: chroma9 = 9'b110110000;
        12'd3367: chroma9 = 9'b110110011;
        12'd3368: chroma9 = 9'b110110110;
        12'd3369: chroma9 = 9'b110111001;
        12'd3370: chroma9 = 9'b110111100;
        12'd3371: chroma9 = 9'b110111111;
        12'd3372: chroma9 = 9'b111000010;
        12'd3373: chroma9 = 9'b111000100;
        12'd3374: chroma9 = 9'b111000110;
        12'd3375: chroma9 = 9'b111001001;
        12'd3376: chroma9 = 9'b111001011;
        12'd3377: chroma9 = 9'b111001101;
        12'd3378: chroma9 = 9'b111001111;
        12'd3379: chroma9 = 9'b111010000;
        12'd3380: chroma9 = 9'b111010010;
        12'd3381: chroma9 = 9'b111010100;
        12'd3382: chroma9 = 9'b111010101;
        12'd3383: chroma9 = 9'b111010110;
        12'd3384: chroma9 = 9'b111010111;
        12'd3385: chroma9 = 9'b111011000;
        12'd3386: chroma9 = 9'b111011001;
        12'd3387: chroma9 = 9'b111011010;
        12'd3388: chroma9 = 9'b111011010;
        12'd3389: chroma9 = 9'b111011011;
        12'd3390: chroma9 = 9'b111011011;
        12'd3391: chroma9 = 9'b111011011;
        12'd3392: chroma9 = 9'b111011011;
        12'd3393: chroma9 = 9'b111011011;
        12'd3394: chroma9 = 9'b111011011;
        12'd3395: chroma9 = 9'b111011011;
        12'd3396: chroma9 = 9'b111011010;
        12'd3397: chroma9 = 9'b111011010;
        12'd3398: chroma9 = 9'b111011001;
        12'd3399: chroma9 = 9'b111011000;
        12'd3400: chroma9 = 9'b111010111;
        12'd3401: chroma9 = 9'b111010110;
        12'd3402: chroma9 = 9'b111010101;
        12'd3403: chroma9 = 9'b111010100;
        12'd3404: chroma9 = 9'b111010010;
        12'd3405: chroma9 = 9'b111010000;
        12'd3406: chroma9 = 9'b111001111;
        12'd3407: chroma9 = 9'b111001101;
        12'd3408: chroma9 = 9'b111001011;
        12'd3409: chroma9 = 9'b111001001;
        12'd3410: chroma9 = 9'b111000110;
        12'd3411: chroma9 = 9'b111000100;
        12'd3412: chroma9 = 9'b111000010;
        12'd3413: chroma9 = 9'b110111111;
        12'd3414: chroma9 = 9'b110111100;
        12'd3415: chroma9 = 9'b110111001;
        12'd3416: chroma9 = 9'b110110110;
        12'd3417: chroma9 = 9'b110110011;
        12'd3418: chroma9 = 9'b110110000;
        12'd3419: chroma9 = 9'b110101101;
        12'd3420: chroma9 = 9'b110101010;
        12'd3421: chroma9 = 9'b110100110;
        12'd3422: chroma9 = 9'b110100011;
        12'd3423: chroma9 = 9'b110011111;
        12'd3424: chroma9 = 9'b110011011;
        12'd3425: chroma9 = 9'b110010111;
        12'd3426: chroma9 = 9'b110010011;
        12'd3427: chroma9 = 9'b110001111;
        12'd3428: chroma9 = 9'b110001011;
        12'd3429: chroma9 = 9'b110000111;
        12'd3430: chroma9 = 9'b110000011;
        12'd3431: chroma9 = 9'b101111110;
        12'd3432: chroma9 = 9'b101111010;
        12'd3433: chroma9 = 9'b101110101;
        12'd3434: chroma9 = 9'b101110001;
        12'd3435: chroma9 = 9'b101101100;
        12'd3436: chroma9 = 9'b101100111;
        12'd3437: chroma9 = 9'b101100010;
        12'd3438: chroma9 = 9'b101011110;
        12'd3439: chroma9 = 9'b101011001;
        12'd3440: chroma9 = 9'b101010100;
        12'd3441: chroma9 = 9'b101001111;
        12'd3442: chroma9 = 9'b101001010;
        12'd3443: chroma9 = 9'b101000101;
        12'd3444: chroma9 = 9'b100111111;
        12'd3445: chroma9 = 9'b100111010;
        12'd3446: chroma9 = 9'b100110101;
        12'd3447: chroma9 = 9'b100110000;
        12'd3448: chroma9 = 9'b100101010;
        12'd3449: chroma9 = 9'b100100101;
        12'd3450: chroma9 = 9'b100100000;
        12'd3451: chroma9 = 9'b100011010;
        12'd3452: chroma9 = 9'b100010101;
        12'd3453: chroma9 = 9'b100010000;
        12'd3454: chroma9 = 9'b100001010;
        12'd3455: chroma9 = 9'b100000101;
        12'd3456: chroma9 = 9'b100000000;
        12'd3457: chroma9 = 9'b011111011;
        12'd3458: chroma9 = 9'b011110110;
        12'd3459: chroma9 = 9'b011110000;
        12'd3460: chroma9 = 9'b011101011;
        12'd3461: chroma9 = 9'b011100110;
        12'd3462: chroma9 = 9'b011100000;
        12'd3463: chroma9 = 9'b011011011;
        12'd3464: chroma9 = 9'b011010110;
        12'd3465: chroma9 = 9'b011010000;
        12'd3466: chroma9 = 9'b011001011;
        12'd3467: chroma9 = 9'b011000110;
        12'd3468: chroma9 = 9'b011000001;
        12'd3469: chroma9 = 9'b010111011;
        12'd3470: chroma9 = 9'b010110110;
        12'd3471: chroma9 = 9'b010110001;
        12'd3472: chroma9 = 9'b010101100;
        12'd3473: chroma9 = 9'b010100111;
        12'd3474: chroma9 = 9'b010100010;
        12'd3475: chroma9 = 9'b010011110;
        12'd3476: chroma9 = 9'b010011001;
        12'd3477: chroma9 = 9'b010010100;
        12'd3478: chroma9 = 9'b010001111;
        12'd3479: chroma9 = 9'b010001011;
        12'd3480: chroma9 = 9'b010000110;
        12'd3481: chroma9 = 9'b010000010;
        12'd3482: chroma9 = 9'b001111101;
        12'd3483: chroma9 = 9'b001111001;
        12'd3484: chroma9 = 9'b001110101;
        12'd3485: chroma9 = 9'b001110001;
        12'd3486: chroma9 = 9'b001101101;
        12'd3487: chroma9 = 9'b001101001;
        12'd3488: chroma9 = 9'b001100101;
        12'd3489: chroma9 = 9'b001100001;
        12'd3490: chroma9 = 9'b001011101;
        12'd3491: chroma9 = 9'b001011010;
        12'd3492: chroma9 = 9'b001010110;
        12'd3493: chroma9 = 9'b001010011;
        12'd3494: chroma9 = 9'b001010000;
        12'd3495: chroma9 = 9'b001001101;
        12'd3496: chroma9 = 9'b001001010;
        12'd3497: chroma9 = 9'b001000111;
        12'd3498: chroma9 = 9'b001000100;
        12'd3499: chroma9 = 9'b001000001;
        12'd3500: chroma9 = 9'b000111110;
        12'd3501: chroma9 = 9'b000111100;
        12'd3502: chroma9 = 9'b000111010;
        12'd3503: chroma9 = 9'b000110111;
        12'd3504: chroma9 = 9'b000110101;
        12'd3505: chroma9 = 9'b000110011;
        12'd3506: chroma9 = 9'b000110001;
        12'd3507: chroma9 = 9'b000110000;
        12'd3508: chroma9 = 9'b000101110;
        12'd3509: chroma9 = 9'b000101100;
        12'd3510: chroma9 = 9'b000101011;
        12'd3511: chroma9 = 9'b000101010;
        12'd3512: chroma9 = 9'b000101001;
        12'd3513: chroma9 = 9'b000101000;
        12'd3514: chroma9 = 9'b000100111;
        12'd3515: chroma9 = 9'b000100110;
        12'd3516: chroma9 = 9'b000100110;
        12'd3517: chroma9 = 9'b000100101;
        12'd3518: chroma9 = 9'b000100101;
        12'd3519: chroma9 = 9'b000100101;
        12'd3520: chroma9 = 9'b000100101;
        12'd3521: chroma9 = 9'b000100101;
        12'd3522: chroma9 = 9'b000100101;
        12'd3523: chroma9 = 9'b000100101;
        12'd3524: chroma9 = 9'b000100110;
        12'd3525: chroma9 = 9'b000100110;
        12'd3526: chroma9 = 9'b000100111;
        12'd3527: chroma9 = 9'b000101000;
        12'd3528: chroma9 = 9'b000101001;
        12'd3529: chroma9 = 9'b000101010;
        12'd3530: chroma9 = 9'b000101011;
        12'd3531: chroma9 = 9'b000101100;
        12'd3532: chroma9 = 9'b000101110;
        12'd3533: chroma9 = 9'b000110000;
        12'd3534: chroma9 = 9'b000110001;
        12'd3535: chroma9 = 9'b000110011;
        12'd3536: chroma9 = 9'b000110101;
        12'd3537: chroma9 = 9'b000110111;
        12'd3538: chroma9 = 9'b000111010;
        12'd3539: chroma9 = 9'b000111100;
        12'd3540: chroma9 = 9'b000111110;
        12'd3541: chroma9 = 9'b001000001;
        12'd3542: chroma9 = 9'b001000100;
        12'd3543: chroma9 = 9'b001000111;
        12'd3544: chroma9 = 9'b001001010;
        12'd3545: chroma9 = 9'b001001101;
        12'd3546: chroma9 = 9'b001010000;
        12'd3547: chroma9 = 9'b001010011;
        12'd3548: chroma9 = 9'b001010110;
        12'd3549: chroma9 = 9'b001011010;
        12'd3550: chroma9 = 9'b001011101;
        12'd3551: chroma9 = 9'b001100001;
        12'd3552: chroma9 = 9'b001100101;
        12'd3553: chroma9 = 9'b001101001;
        12'd3554: chroma9 = 9'b001101101;
        12'd3555: chroma9 = 9'b001110001;
        12'd3556: chroma9 = 9'b001110101;
        12'd3557: chroma9 = 9'b001111001;
        12'd3558: chroma9 = 9'b001111101;
        12'd3559: chroma9 = 9'b010000010;
        12'd3560: chroma9 = 9'b010000110;
        12'd3561: chroma9 = 9'b010001011;
        12'd3562: chroma9 = 9'b010001111;
        12'd3563: chroma9 = 9'b010010100;
        12'd3564: chroma9 = 9'b010011001;
        12'd3565: chroma9 = 9'b010011110;
        12'd3566: chroma9 = 9'b010100010;
        12'd3567: chroma9 = 9'b010100111;
        12'd3568: chroma9 = 9'b010101100;
        12'd3569: chroma9 = 9'b010110001;
        12'd3570: chroma9 = 9'b010110110;
        12'd3571: chroma9 = 9'b010111011;
        12'd3572: chroma9 = 9'b011000001;
        12'd3573: chroma9 = 9'b011000110;
        12'd3574: chroma9 = 9'b011001011;
        12'd3575: chroma9 = 9'b011010000;
        12'd3576: chroma9 = 9'b011010110;
        12'd3577: chroma9 = 9'b011011011;
        12'd3578: chroma9 = 9'b011100000;
        12'd3579: chroma9 = 9'b011100110;
        12'd3580: chroma9 = 9'b011101011;
        12'd3581: chroma9 = 9'b011110000;
        12'd3582: chroma9 = 9'b011110110;
        12'd3583: chroma9 = 9'b011111011;
        12'd3584: chroma9 = 9'b100000000;
        12'd3585: chroma9 = 9'b100000101;
        12'd3586: chroma9 = 9'b100001011;
        12'd3587: chroma9 = 9'b100010001;
        12'd3588: chroma9 = 9'b100010111;
        12'd3589: chroma9 = 9'b100011100;
        12'd3590: chroma9 = 9'b100100010;
        12'd3591: chroma9 = 9'b100101000;
        12'd3592: chroma9 = 9'b100101101;
        12'd3593: chroma9 = 9'b100110011;
        12'd3594: chroma9 = 9'b100111001;
        12'd3595: chroma9 = 9'b100111110;
        12'd3596: chroma9 = 9'b101000100;
        12'd3597: chroma9 = 9'b101001001;
        12'd3598: chroma9 = 9'b101001111;
        12'd3599: chroma9 = 9'b101010100;
        12'd3600: chroma9 = 9'b101011001;
        12'd3601: chroma9 = 9'b101011111;
        12'd3602: chroma9 = 9'b101100100;
        12'd3603: chroma9 = 9'b101101001;
        12'd3604: chroma9 = 9'b101101110;
        12'd3605: chroma9 = 9'b101110011;
        12'd3606: chroma9 = 9'b101111000;
        12'd3607: chroma9 = 9'b101111101;
        12'd3608: chroma9 = 9'b110000010;
        12'd3609: chroma9 = 9'b110000111;
        12'd3610: chroma9 = 9'b110001011;
        12'd3611: chroma9 = 9'b110010000;
        12'd3612: chroma9 = 9'b110010101;
        12'd3613: chroma9 = 9'b110011001;
        12'd3614: chroma9 = 9'b110011101;
        12'd3615: chroma9 = 9'b110100010;
        12'd3616: chroma9 = 9'b110100110;
        12'd3617: chroma9 = 9'b110101010;
        12'd3618: chroma9 = 9'b110101110;
        12'd3619: chroma9 = 9'b110110001;
        12'd3620: chroma9 = 9'b110110101;
        12'd3621: chroma9 = 9'b110111001;
        12'd3622: chroma9 = 9'b110111100;
        12'd3623: chroma9 = 9'b111000000;
        12'd3624: chroma9 = 9'b111000011;
        12'd3625: chroma9 = 9'b111000110;
        12'd3626: chroma9 = 9'b111001001;
        12'd3627: chroma9 = 9'b111001100;
        12'd3628: chroma9 = 9'b111001111;
        12'd3629: chroma9 = 9'b111010001;
        12'd3630: chroma9 = 9'b111010100;
        12'd3631: chroma9 = 9'b111010110;
        12'd3632: chroma9 = 9'b111011001;
        12'd3633: chroma9 = 9'b111011011;
        12'd3634: chroma9 = 9'b111011101;
        12'd3635: chroma9 = 9'b111011111;
        12'd3636: chroma9 = 9'b111100000;
        12'd3637: chroma9 = 9'b111100010;
        12'd3638: chroma9 = 9'b111100011;
        12'd3639: chroma9 = 9'b111100101;
        12'd3640: chroma9 = 9'b111100110;
        12'd3641: chroma9 = 9'b111100111;
        12'd3642: chroma9 = 9'b111101000;
        12'd3643: chroma9 = 9'b111101001;
        12'd3644: chroma9 = 9'b111101001;
        12'd3645: chroma9 = 9'b111101010;
        12'd3646: chroma9 = 9'b111101010;
        12'd3647: chroma9 = 9'b111101010;
        12'd3648: chroma9 = 9'b111101010;
        12'd3649: chroma9 = 9'b111101010;
        12'd3650: chroma9 = 9'b111101010;
        12'd3651: chroma9 = 9'b111101010;
        12'd3652: chroma9 = 9'b111101001;
        12'd3653: chroma9 = 9'b111101001;
        12'd3654: chroma9 = 9'b111101000;
        12'd3655: chroma9 = 9'b111100111;
        12'd3656: chroma9 = 9'b111100110;
        12'd3657: chroma9 = 9'b111100101;
        12'd3658: chroma9 = 9'b111100011;
        12'd3659: chroma9 = 9'b111100010;
        12'd3660: chroma9 = 9'b111100000;
        12'd3661: chroma9 = 9'b111011111;
        12'd3662: chroma9 = 9'b111011101;
        12'd3663: chroma9 = 9'b111011011;
        12'd3664: chroma9 = 9'b111011001;
        12'd3665: chroma9 = 9'b111010110;
        12'd3666: chroma9 = 9'b111010100;
        12'd3667: chroma9 = 9'b111010001;
        12'd3668: chroma9 = 9'b111001111;
        12'd3669: chroma9 = 9'b111001100;
        12'd3670: chroma9 = 9'b111001001;
        12'd3671: chroma9 = 9'b111000110;
        12'd3672: chroma9 = 9'b111000011;
        12'd3673: chroma9 = 9'b111000000;
        12'd3674: chroma9 = 9'b110111100;
        12'd3675: chroma9 = 9'b110111001;
        12'd3676: chroma9 = 9'b110110101;
        12'd3677: chroma9 = 9'b110110001;
        12'd3678: chroma9 = 9'b110101110;
        12'd3679: chroma9 = 9'b110101010;
        12'd3680: chroma9 = 9'b110100110;
        12'd3681: chroma9 = 9'b110100010;
        12'd3682: chroma9 = 9'b110011101;
        12'd3683: chroma9 = 9'b110011001;
        12'd3684: chroma9 = 9'b110010101;
        12'd3685: chroma9 = 9'b110010000;
        12'd3686: chroma9 = 9'b110001011;
        12'd3687: chroma9 = 9'b110000111;
        12'd3688: chroma9 = 9'b110000010;
        12'd3689: chroma9 = 9'b101111101;
        12'd3690: chroma9 = 9'b101111000;
        12'd3691: chroma9 = 9'b101110011;
        12'd3692: chroma9 = 9'b101101110;
        12'd3693: chroma9 = 9'b101101001;
        12'd3694: chroma9 = 9'b101100100;
        12'd3695: chroma9 = 9'b101011111;
        12'd3696: chroma9 = 9'b101011001;
        12'd3697: chroma9 = 9'b101010100;
        12'd3698: chroma9 = 9'b101001111;
        12'd3699: chroma9 = 9'b101001001;
        12'd3700: chroma9 = 9'b101000100;
        12'd3701: chroma9 = 9'b100111110;
        12'd3702: chroma9 = 9'b100111001;
        12'd3703: chroma9 = 9'b100110011;
        12'd3704: chroma9 = 9'b100101101;
        12'd3705: chroma9 = 9'b100101000;
        12'd3706: chroma9 = 9'b100100010;
        12'd3707: chroma9 = 9'b100011100;
        12'd3708: chroma9 = 9'b100010111;
        12'd3709: chroma9 = 9'b100010001;
        12'd3710: chroma9 = 9'b100001011;
        12'd3711: chroma9 = 9'b100000101;
        12'd3712: chroma9 = 9'b100000000;
        12'd3713: chroma9 = 9'b011111011;
        12'd3714: chroma9 = 9'b011110101;
        12'd3715: chroma9 = 9'b011101111;
        12'd3716: chroma9 = 9'b011101001;
        12'd3717: chroma9 = 9'b011100100;
        12'd3718: chroma9 = 9'b011011110;
        12'd3719: chroma9 = 9'b011011000;
        12'd3720: chroma9 = 9'b011010011;
        12'd3721: chroma9 = 9'b011001101;
        12'd3722: chroma9 = 9'b011000111;
        12'd3723: chroma9 = 9'b011000010;
        12'd3724: chroma9 = 9'b010111100;
        12'd3725: chroma9 = 9'b010110111;
        12'd3726: chroma9 = 9'b010110001;
        12'd3727: chroma9 = 9'b010101100;
        12'd3728: chroma9 = 9'b010100111;
        12'd3729: chroma9 = 9'b010100001;
        12'd3730: chroma9 = 9'b010011100;
        12'd3731: chroma9 = 9'b010010111;
        12'd3732: chroma9 = 9'b010010010;
        12'd3733: chroma9 = 9'b010001101;
        12'd3734: chroma9 = 9'b010001000;
        12'd3735: chroma9 = 9'b010000011;
        12'd3736: chroma9 = 9'b001111110;
        12'd3737: chroma9 = 9'b001111001;
        12'd3738: chroma9 = 9'b001110101;
        12'd3739: chroma9 = 9'b001110000;
        12'd3740: chroma9 = 9'b001101011;
        12'd3741: chroma9 = 9'b001100111;
        12'd3742: chroma9 = 9'b001100011;
        12'd3743: chroma9 = 9'b001011110;
        12'd3744: chroma9 = 9'b001011010;
        12'd3745: chroma9 = 9'b001010110;
        12'd3746: chroma9 = 9'b001010010;
        12'd3747: chroma9 = 9'b001001111;
        12'd3748: chroma9 = 9'b001001011;
        12'd3749: chroma9 = 9'b001000111;
        12'd3750: chroma9 = 9'b001000100;
        12'd3751: chroma9 = 9'b001000000;
        12'd3752: chroma9 = 9'b000111101;
        12'd3753: chroma9 = 9'b000111010;
        12'd3754: chroma9 = 9'b000110111;
        12'd3755: chroma9 = 9'b000110100;
        12'd3756: chroma9 = 9'b000110001;
        12'd3757: chroma9 = 9'b000101111;
        12'd3758: chroma9 = 9'b000101100;
        12'd3759: chroma9 = 9'b000101010;
        12'd3760: chroma9 = 9'b000100111;
        12'd3761: chroma9 = 9'b000100101;
        12'd3762: chroma9 = 9'b000100011;
        12'd3763: chroma9 = 9'b000100001;
        12'd3764: chroma9 = 9'b000100000;
        12'd3765: chroma9 = 9'b000011110;
        12'd3766: chroma9 = 9'b000011101;
        12'd3767: chroma9 = 9'b000011011;
        12'd3768: chroma9 = 9'b000011010;
        12'd3769: chroma9 = 9'b000011001;
        12'd3770: chroma9 = 9'b000011000;
        12'd3771: chroma9 = 9'b000010111;
        12'd3772: chroma9 = 9'b000010111;
        12'd3773: chroma9 = 9'b000010110;
        12'd3774: chroma9 = 9'b000010110;
        12'd3775: chroma9 = 9'b000010110;
        12'd3776: chroma9 = 9'b000010110;
        12'd3777: chroma9 = 9'b000010110;
        12'd3778: chroma9 = 9'b000010110;
        12'd3779: chroma9 = 9'b000010110;
        12'd3780: chroma9 = 9'b000010111;
        12'd3781: chroma9 = 9'b000010111;
        12'd3782: chroma9 = 9'b000011000;
        12'd3783: chroma9 = 9'b000011001;
        12'd3784: chroma9 = 9'b000011010;
        12'd3785: chroma9 = 9'b000011011;
        12'd3786: chroma9 = 9'b000011101;
        12'd3787: chroma9 = 9'b000011110;
        12'd3788: chroma9 = 9'b000100000;
        12'd3789: chroma9 = 9'b000100001;
        12'd3790: chroma9 = 9'b000100011;
        12'd3791: chroma9 = 9'b000100101;
        12'd3792: chroma9 = 9'b000100111;
        12'd3793: chroma9 = 9'b000101010;
        12'd3794: chroma9 = 9'b000101100;
        12'd3795: chroma9 = 9'b000101111;
        12'd3796: chroma9 = 9'b000110001;
        12'd3797: chroma9 = 9'b000110100;
        12'd3798: chroma9 = 9'b000110111;
        12'd3799: chroma9 = 9'b000111010;
        12'd3800: chroma9 = 9'b000111101;
        12'd3801: chroma9 = 9'b001000000;
        12'd3802: chroma9 = 9'b001000100;
        12'd3803: chroma9 = 9'b001000111;
        12'd3804: chroma9 = 9'b001001011;
        12'd3805: chroma9 = 9'b001001111;
        12'd3806: chroma9 = 9'b001010010;
        12'd3807: chroma9 = 9'b001010110;
        12'd3808: chroma9 = 9'b001011010;
        12'd3809: chroma9 = 9'b001011110;
        12'd3810: chroma9 = 9'b001100011;
        12'd3811: chroma9 = 9'b001100111;
        12'd3812: chroma9 = 9'b001101011;
        12'd3813: chroma9 = 9'b001110000;
        12'd3814: chroma9 = 9'b001110101;
        12'd3815: chroma9 = 9'b001111001;
        12'd3816: chroma9 = 9'b001111110;
        12'd3817: chroma9 = 9'b010000011;
        12'd3818: chroma9 = 9'b010001000;
        12'd3819: chroma9 = 9'b010001101;
        12'd3820: chroma9 = 9'b010010010;
        12'd3821: chroma9 = 9'b010010111;
        12'd3822: chroma9 = 9'b010011100;
        12'd3823: chroma9 = 9'b010100001;
        12'd3824: chroma9 = 9'b010100111;
        12'd3825: chroma9 = 9'b010101100;
        12'd3826: chroma9 = 9'b010110001;
        12'd3827: chroma9 = 9'b010110111;
        12'd3828: chroma9 = 9'b010111100;
        12'd3829: chroma9 = 9'b011000010;
        12'd3830: chroma9 = 9'b011000111;
        12'd3831: chroma9 = 9'b011001101;
        12'd3832: chroma9 = 9'b011010011;
        12'd3833: chroma9 = 9'b011011000;
        12'd3834: chroma9 = 9'b011011110;
        12'd3835: chroma9 = 9'b011100100;
        12'd3836: chroma9 = 9'b011101001;
        12'd3837: chroma9 = 9'b011101111;
        12'd3838: chroma9 = 9'b011110101;
        12'd3839: chroma9 = 9'b011111011;
        12'd3840: chroma9 = 9'b100000000;
        12'd3841: chroma9 = 9'b100000110;
        12'd3842: chroma9 = 9'b100001100;
        12'd3843: chroma9 = 9'b100010010;
        12'd3844: chroma9 = 9'b100011000;
        12'd3845: chroma9 = 9'b100011110;
        12'd3846: chroma9 = 9'b100100100;
        12'd3847: chroma9 = 9'b100101010;
        12'd3848: chroma9 = 9'b100110000;
        12'd3849: chroma9 = 9'b100110110;
        12'd3850: chroma9 = 9'b100111100;
        12'd3851: chroma9 = 9'b101000010;
        12'd3852: chroma9 = 9'b101001000;
        12'd3853: chroma9 = 9'b101001110;
        12'd3854: chroma9 = 9'b101010100;
        12'd3855: chroma9 = 9'b101011001;
        12'd3856: chroma9 = 9'b101011111;
        12'd3857: chroma9 = 9'b101100101;
        12'd3858: chroma9 = 9'b101101010;
        12'd3859: chroma9 = 9'b101110000;
        12'd3860: chroma9 = 9'b101110101;
        12'd3861: chroma9 = 9'b101111011;
        12'd3862: chroma9 = 9'b110000000;
        12'd3863: chroma9 = 9'b110000101;
        12'd3864: chroma9 = 9'b110001010;
        12'd3865: chroma9 = 9'b110001111;
        12'd3866: chroma9 = 9'b110010100;
        12'd3867: chroma9 = 9'b110011001;
        12'd3868: chroma9 = 9'b110011110;
        12'd3869: chroma9 = 9'b110100011;
        12'd3870: chroma9 = 9'b110100111;
        12'd3871: chroma9 = 9'b110101100;
        12'd3872: chroma9 = 9'b110110000;
        12'd3873: chroma9 = 9'b110110101;
        12'd3874: chroma9 = 9'b110111001;
        12'd3875: chroma9 = 9'b110111101;
        12'd3876: chroma9 = 9'b111000001;
        12'd3877: chroma9 = 9'b111000101;
        12'd3878: chroma9 = 9'b111001000;
        12'd3879: chroma9 = 9'b111001100;
        12'd3880: chroma9 = 9'b111001111;
        12'd3881: chroma9 = 9'b111010011;
        12'd3882: chroma9 = 9'b111010110;
        12'd3883: chroma9 = 9'b111011001;
        12'd3884: chroma9 = 9'b111011100;
        12'd3885: chroma9 = 9'b111011111;
        12'd3886: chroma9 = 9'b111100001;
        12'd3887: chroma9 = 9'b111100100;
        12'd3888: chroma9 = 9'b111100110;
        12'd3889: chroma9 = 9'b111101001;
        12'd3890: chroma9 = 9'b111101011;
        12'd3891: chroma9 = 9'b111101101;
        12'd3892: chroma9 = 9'b111101111;
        12'd3893: chroma9 = 9'b111110000;
        12'd3894: chroma9 = 9'b111110010;
        12'd3895: chroma9 = 9'b111110011;
        12'd3896: chroma9 = 9'b111110101;
        12'd3897: chroma9 = 9'b111110110;
        12'd3898: chroma9 = 9'b111110111;
        12'd3899: chroma9 = 9'b111111000;
        12'd3900: chroma9 = 9'b111111000;
        12'd3901: chroma9 = 9'b111111001;
        12'd3902: chroma9 = 9'b111111001;
        12'd3903: chroma9 = 9'b111111001;
        12'd3904: chroma9 = 9'b111111001;
        12'd3905: chroma9 = 9'b111111001;
        12'd3906: chroma9 = 9'b111111001;
        12'd3907: chroma9 = 9'b111111001;
        12'd3908: chroma9 = 9'b111111000;
        12'd3909: chroma9 = 9'b111111000;
        12'd3910: chroma9 = 9'b111110111;
        12'd3911: chroma9 = 9'b111110110;
        12'd3912: chroma9 = 9'b111110101;
        12'd3913: chroma9 = 9'b111110011;
        12'd3914: chroma9 = 9'b111110010;
        12'd3915: chroma9 = 9'b111110000;
        12'd3916: chroma9 = 9'b111101111;
        12'd3917: chroma9 = 9'b111101101;
        12'd3918: chroma9 = 9'b111101011;
        12'd3919: chroma9 = 9'b111101001;
        12'd3920: chroma9 = 9'b111100110;
        12'd3921: chroma9 = 9'b111100100;
        12'd3922: chroma9 = 9'b111100001;
        12'd3923: chroma9 = 9'b111011111;
        12'd3924: chroma9 = 9'b111011100;
        12'd3925: chroma9 = 9'b111011001;
        12'd3926: chroma9 = 9'b111010110;
        12'd3927: chroma9 = 9'b111010011;
        12'd3928: chroma9 = 9'b111001111;
        12'd3929: chroma9 = 9'b111001100;
        12'd3930: chroma9 = 9'b111001000;
        12'd3931: chroma9 = 9'b111000101;
        12'd3932: chroma9 = 9'b111000001;
        12'd3933: chroma9 = 9'b110111101;
        12'd3934: chroma9 = 9'b110111001;
        12'd3935: chroma9 = 9'b110110101;
        12'd3936: chroma9 = 9'b110110000;
        12'd3937: chroma9 = 9'b110101100;
        12'd3938: chroma9 = 9'b110100111;
        12'd3939: chroma9 = 9'b110100011;
        12'd3940: chroma9 = 9'b110011110;
        12'd3941: chroma9 = 9'b110011001;
        12'd3942: chroma9 = 9'b110010100;
        12'd3943: chroma9 = 9'b110001111;
        12'd3944: chroma9 = 9'b110001010;
        12'd3945: chroma9 = 9'b110000101;
        12'd3946: chroma9 = 9'b110000000;
        12'd3947: chroma9 = 9'b101111011;
        12'd3948: chroma9 = 9'b101110101;
        12'd3949: chroma9 = 9'b101110000;
        12'd3950: chroma9 = 9'b101101010;
        12'd3951: chroma9 = 9'b101100101;
        12'd3952: chroma9 = 9'b101011111;
        12'd3953: chroma9 = 9'b101011001;
        12'd3954: chroma9 = 9'b101010100;
        12'd3955: chroma9 = 9'b101001110;
        12'd3956: chroma9 = 9'b101001000;
        12'd3957: chroma9 = 9'b101000010;
        12'd3958: chroma9 = 9'b100111100;
        12'd3959: chroma9 = 9'b100110110;
        12'd3960: chroma9 = 9'b100110000;
        12'd3961: chroma9 = 9'b100101010;
        12'd3962: chroma9 = 9'b100100100;
        12'd3963: chroma9 = 9'b100011110;
        12'd3964: chroma9 = 9'b100011000;
        12'd3965: chroma9 = 9'b100010010;
        12'd3966: chroma9 = 9'b100001100;
        12'd3967: chroma9 = 9'b100000110;
        12'd3968: chroma9 = 9'b100000000;
        12'd3969: chroma9 = 9'b011111010;
        12'd3970: chroma9 = 9'b011110100;
        12'd3971: chroma9 = 9'b011101110;
        12'd3972: chroma9 = 9'b011101000;
        12'd3973: chroma9 = 9'b011100010;
        12'd3974: chroma9 = 9'b011011100;
        12'd3975: chroma9 = 9'b011010110;
        12'd3976: chroma9 = 9'b011010000;
        12'd3977: chroma9 = 9'b011001010;
        12'd3978: chroma9 = 9'b011000100;
        12'd3979: chroma9 = 9'b010111110;
        12'd3980: chroma9 = 9'b010111000;
        12'd3981: chroma9 = 9'b010110010;
        12'd3982: chroma9 = 9'b010101100;
        12'd3983: chroma9 = 9'b010100111;
        12'd3984: chroma9 = 9'b010100001;
        12'd3985: chroma9 = 9'b010011011;
        12'd3986: chroma9 = 9'b010010110;
        12'd3987: chroma9 = 9'b010010000;
        12'd3988: chroma9 = 9'b010001011;
        12'd3989: chroma9 = 9'b010000101;
        12'd3990: chroma9 = 9'b010000000;
        12'd3991: chroma9 = 9'b001111011;
        12'd3992: chroma9 = 9'b001110110;
        12'd3993: chroma9 = 9'b001110001;
        12'd3994: chroma9 = 9'b001101100;
        12'd3995: chroma9 = 9'b001100111;
        12'd3996: chroma9 = 9'b001100010;
        12'd3997: chroma9 = 9'b001011101;
        12'd3998: chroma9 = 9'b001011001;
        12'd3999: chroma9 = 9'b001010100;
        12'd4000: chroma9 = 9'b001010000;
        12'd4001: chroma9 = 9'b001001011;
        12'd4002: chroma9 = 9'b001000111;
        12'd4003: chroma9 = 9'b001000011;
        12'd4004: chroma9 = 9'b000111111;
        12'd4005: chroma9 = 9'b000111011;
        12'd4006: chroma9 = 9'b000111000;
        12'd4007: chroma9 = 9'b000110100;
        12'd4008: chroma9 = 9'b000110001;
        12'd4009: chroma9 = 9'b000101101;
        12'd4010: chroma9 = 9'b000101010;
        12'd4011: chroma9 = 9'b000100111;
        12'd4012: chroma9 = 9'b000100100;
        12'd4013: chroma9 = 9'b000100001;
        12'd4014: chroma9 = 9'b000011111;
        12'd4015: chroma9 = 9'b000011100;
        12'd4016: chroma9 = 9'b000011010;
        12'd4017: chroma9 = 9'b000010111;
        12'd4018: chroma9 = 9'b000010101;
        12'd4019: chroma9 = 9'b000010011;
        12'd4020: chroma9 = 9'b000010001;
        12'd4021: chroma9 = 9'b000010000;
        12'd4022: chroma9 = 9'b000001110;
        12'd4023: chroma9 = 9'b000001101;
        12'd4024: chroma9 = 9'b000001011;
        12'd4025: chroma9 = 9'b000001010;
        12'd4026: chroma9 = 9'b000001001;
        12'd4027: chroma9 = 9'b000001000;
        12'd4028: chroma9 = 9'b000001000;
        12'd4029: chroma9 = 9'b000000111;
        12'd4030: chroma9 = 9'b000000111;
        12'd4031: chroma9 = 9'b000000111;
        12'd4032: chroma9 = 9'b000000111;
        12'd4033: chroma9 = 9'b000000111;
        12'd4034: chroma9 = 9'b000000111;
        12'd4035: chroma9 = 9'b000000111;
        12'd4036: chroma9 = 9'b000001000;
        12'd4037: chroma9 = 9'b000001000;
        12'd4038: chroma9 = 9'b000001001;
        12'd4039: chroma9 = 9'b000001010;
        12'd4040: chroma9 = 9'b000001011;
        12'd4041: chroma9 = 9'b000001101;
        12'd4042: chroma9 = 9'b000001110;
        12'd4043: chroma9 = 9'b000010000;
        12'd4044: chroma9 = 9'b000010001;
        12'd4045: chroma9 = 9'b000010011;
        12'd4046: chroma9 = 9'b000010101;
        12'd4047: chroma9 = 9'b000010111;
        12'd4048: chroma9 = 9'b000011010;
        12'd4049: chroma9 = 9'b000011100;
        12'd4050: chroma9 = 9'b000011111;
        12'd4051: chroma9 = 9'b000100001;
        12'd4052: chroma9 = 9'b000100100;
        12'd4053: chroma9 = 9'b000100111;
        12'd4054: chroma9 = 9'b000101010;
        12'd4055: chroma9 = 9'b000101101;
        12'd4056: chroma9 = 9'b000110001;
        12'd4057: chroma9 = 9'b000110100;
        12'd4058: chroma9 = 9'b000111000;
        12'd4059: chroma9 = 9'b000111011;
        12'd4060: chroma9 = 9'b000111111;
        12'd4061: chroma9 = 9'b001000011;
        12'd4062: chroma9 = 9'b001000111;
        12'd4063: chroma9 = 9'b001001011;
        12'd4064: chroma9 = 9'b001010000;
        12'd4065: chroma9 = 9'b001010100;
        12'd4066: chroma9 = 9'b001011001;
        12'd4067: chroma9 = 9'b001011101;
        12'd4068: chroma9 = 9'b001100010;
        12'd4069: chroma9 = 9'b001100111;
        12'd4070: chroma9 = 9'b001101100;
        12'd4071: chroma9 = 9'b001110001;
        12'd4072: chroma9 = 9'b001110110;
        12'd4073: chroma9 = 9'b001111011;
        12'd4074: chroma9 = 9'b010000000;
        12'd4075: chroma9 = 9'b010000101;
        12'd4076: chroma9 = 9'b010001011;
        12'd4077: chroma9 = 9'b010010000;
        12'd4078: chroma9 = 9'b010010110;
        12'd4079: chroma9 = 9'b010011011;
        12'd4080: chroma9 = 9'b010100001;
        12'd4081: chroma9 = 9'b010100111;
        12'd4082: chroma9 = 9'b010101100;
        12'd4083: chroma9 = 9'b010110010;
        12'd4084: chroma9 = 9'b010111000;
        12'd4085: chroma9 = 9'b010111110;
        12'd4086: chroma9 = 9'b011000100;
        12'd4087: chroma9 = 9'b011001010;
        12'd4088: chroma9 = 9'b011010000;
        12'd4089: chroma9 = 9'b011010110;
        12'd4090: chroma9 = 9'b011011100;
        12'd4091: chroma9 = 9'b011100010;
        12'd4092: chroma9 = 9'b011101000;
        12'd4093: chroma9 = 9'b011101110;
        12'd4094: chroma9 = 9'b011110100;
        12'd4095: chroma9 = 9'b011111010;
    endcase
end
`endif

endmodule
