`ifndef config_vh_
`define config_vh_

`define VERSION_MAJOR 8'd1
`define VERSION_MINOR 8'd5

`define EFINIX
`define VARIANT_SUFFIX_1 8'd76
`define VARIANT_SUFFIX_2 8'd72
`define VARIANT_SUFFIX_3 8'd0
`define VARIANT_SUFFIX_4 8'd0
`define WITH_EXTENSIONS 1
`define GEN_LUMA_CHROMA 1
`define CONFIGURABLE_RGB 1
`define CONFIGURABLE_LUMAS 1
`define HIRES_MODES 1
`define WITH_MATH 1
`define WITH_RAM 1
`define WITH_64K 1
`define HAVE_EEPROM 1
`define HAVE_FLASH 1
`define WITH_BLITTER 1

`endif // config_vh_
