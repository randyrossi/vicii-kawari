// Init sequence code for board with MCU.
// In this config, we use the MCU's EEPROM
// to store/retrieve settings. For chip, the MCU
// is simply setting the incoming chip_ext lines
// hi/lo depending on what chip was persisted
// in EEPROM (on MCU). We just hold reset for a
// while and then switch chip half way through.
//
// All other settings are sent via serial link
// after cclk goes high (indicating loading
// is complete by MCU) and are handled in
// registers_ram.v

`ifndef SIMULATOR_BOARD
// @ 14Mhz, 1/14000000*2^21 = ~ 149ms
`define RESET_CTR_TOP_BIT 20
`define RESET_CTR_INC 21'd1
`define RESET_LATCH_POINT 21'b010000000000000000000
`else
// For simluator, have a much shorter reset period 
`define RESET_CTR_TOP_BIT 7
`define RESET_CTR_INC 7'd1
`define RESET_LATCH_POINT 8'b01000000
`endif

reg [`RESET_CTR_TOP_BIT:0] rstcntr = 0;
wire internal_rst = !rstcntr[`RESET_CTR_TOP_BIT];

always @(posedge clk_dot4x)
begin
    if (internal_rst)
        rstcntr <= rstcntr + `RESET_CTR_INC;
    if (rstcntr == `RESET_LATCH_POINT) begin
        $display("chip <= %d", chip_ext);
        chip <= chip_ext;
    end
end

// Take design out of reset when internal_rst is high
always @(posedge clk_dot4x) rst <= internal_rst;
