`ifndef common_vh_
`define common_vh_

typedef enum [1:0] { CHIP6567R8, CHIP6567R56A, CHIP6569, CHIPUNUSED} chip_type;

`define TRUE	1'b1
`define FALSE	1'b0

`endif // common_vh_